
module FullAdder_0 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2017 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2018 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2019 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2020 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2021 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2022 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2023 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2024 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2025 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2026 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2027 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2028 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2029 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2030 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2031 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2032 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2033 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2034 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2035 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2036 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2037 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2038 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2039 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2040 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2041 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2042 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2043 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2044 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2045 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2046 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2047 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_0 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_0 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_2047 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_2046 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_2045 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_2044 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_2043 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_2042 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_2041 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_2040 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_2039 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_2038 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_2037 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_2036 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_2035 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_2034 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_2033 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_2032 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_2031 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_2030 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_2029 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_2028 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_2027 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_2026 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_2025 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_2024 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_2023 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_2022 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_2021 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_2020 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_2019 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_2018 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_2017 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1985 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1986 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1987 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1988 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1989 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1990 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1991 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1992 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1993 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1994 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1995 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1996 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1997 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1998 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1999 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2000 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2001 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2002 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2003 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2004 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2005 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2006 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2007 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2008 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2009 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2010 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2011 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2012 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2013 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2014 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2015 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2016 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_63 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_2016 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_2015 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_2014 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_2013 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_2012 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_2011 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_2010 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_2009 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_2008 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_2007 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_2006 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_2005 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_2004 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_2003 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_2002 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_2001 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_2000 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1999 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1998 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1997 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1996 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1995 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1994 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1993 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1992 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1991 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1990 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1989 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1988 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1987 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1986 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1985 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_0 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n65, n66, n67, n68;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_0 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_63 sub ( .a(a), .b({n33, n34, n35, n36, n37, n38, n39, n40, n41, 
        n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, 
        n56, n57, n58, n59, n60, n61, n62, n63, n64}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n64) );
  INV_X1 U72 ( .A(m[1]), .ZN(n63) );
  INV_X1 U73 ( .A(m[2]), .ZN(n62) );
  INV_X1 U74 ( .A(m[3]), .ZN(n61) );
  INV_X1 U75 ( .A(m[4]), .ZN(n60) );
  INV_X1 U76 ( .A(m[5]), .ZN(n59) );
  INV_X1 U77 ( .A(m[6]), .ZN(n58) );
  INV_X1 U78 ( .A(m[7]), .ZN(n57) );
  INV_X1 U79 ( .A(m[8]), .ZN(n56) );
  INV_X1 U80 ( .A(m[9]), .ZN(n55) );
  INV_X1 U81 ( .A(m[10]), .ZN(n54) );
  INV_X1 U82 ( .A(m[11]), .ZN(n53) );
  INV_X1 U83 ( .A(m[12]), .ZN(n52) );
  INV_X1 U84 ( .A(m[13]), .ZN(n51) );
  INV_X1 U85 ( .A(m[14]), .ZN(n50) );
  INV_X1 U86 ( .A(m[15]), .ZN(n49) );
  INV_X1 U87 ( .A(m[16]), .ZN(n48) );
  INV_X1 U88 ( .A(m[17]), .ZN(n47) );
  INV_X1 U89 ( .A(m[18]), .ZN(n46) );
  INV_X1 U90 ( .A(m[19]), .ZN(n45) );
  INV_X1 U91 ( .A(m[20]), .ZN(n44) );
  INV_X1 U92 ( .A(m[21]), .ZN(n43) );
  INV_X1 U93 ( .A(m[22]), .ZN(n42) );
  INV_X1 U94 ( .A(m[23]), .ZN(n41) );
  INV_X1 U95 ( .A(m[24]), .ZN(n40) );
  INV_X1 U96 ( .A(m[25]), .ZN(n39) );
  INV_X1 U97 ( .A(m[26]), .ZN(n38) );
  INV_X1 U98 ( .A(m[27]), .ZN(n37) );
  INV_X1 U99 ( .A(m[28]), .ZN(n36) );
  INV_X1 U100 ( .A(m[29]), .ZN(n35) );
  INV_X1 U101 ( .A(m[30]), .ZN(n34) );
  INV_X1 U102 ( .A(m[31]), .ZN(n33) );
endmodule


module FullAdder_1 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_3 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_4 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_5 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_6 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_7 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_8 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_9 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_10 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_11 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_12 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_13 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_14 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_15 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_16 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_17 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_18 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_19 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_20 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_21 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_22 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_23 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_24 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_25 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_26 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_27 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_28 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_29 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_30 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_31 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_32 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_1 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_32 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_31 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_30 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_29 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_28 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_27 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_26 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_25 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_24 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_23 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_22 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_21 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_20 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_19 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_18 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_17 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_16 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_15 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_14 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_13 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_12 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_11 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_10 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_9 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_8 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_7 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_6 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_5 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_4 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_3 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_2 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), 
        .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_33 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_34 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_35 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_36 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_37 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_38 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_39 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_40 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_41 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_42 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_43 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_44 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_45 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_46 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_47 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_48 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_49 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_50 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_51 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_52 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_53 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_54 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_55 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_56 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_57 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_58 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_59 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_60 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_61 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_62 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_63 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_64 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_2 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_64 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_63 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_62 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_61 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_60 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_59 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_58 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_57 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_56 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_55 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_54 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_53 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_52 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_51 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_50 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_49 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_48 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_47 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_46 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_45 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_44 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_43 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_42 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_41 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_40 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_39 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_38 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_37 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_36 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_35 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_34 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_33 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), 
        .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_1 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_2 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_1 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_65 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_66 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_67 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_68 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_69 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_70 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_71 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_72 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_73 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_74 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_75 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_76 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_77 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_78 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_79 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_80 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_81 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_82 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_83 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_84 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_85 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_86 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_87 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_88 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_89 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_90 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_91 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_92 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_93 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_94 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_95 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_96 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_3 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_96 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_95 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_94 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_93 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_92 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_91 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_90 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_89 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_88 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_87 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_86 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_85 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_84 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_83 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_82 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_81 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_80 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_79 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_78 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_77 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_76 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_75 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_74 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_73 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_72 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_71 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_70 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_69 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_68 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_67 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_66 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_65 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), 
        .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_97 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_98 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_99 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_100 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_101 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_102 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_103 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_104 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_105 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_106 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_107 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_108 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_109 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_110 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_111 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_112 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_113 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_114 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_115 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_116 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_117 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_118 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_119 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_120 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_121 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_122 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_123 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_124 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_125 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_126 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_127 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_128 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_4 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_128 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_127 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_126 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_125 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_124 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_123 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_122 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_121 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_120 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_119 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_118 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_117 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_116 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_115 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_114 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_113 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_112 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_111 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_110 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_109 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_108 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_107 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_106 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_105 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_104 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_103 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_102 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_101 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_100 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_99 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_98 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_97 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), 
        .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_2 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_4 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_3 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_129 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_130 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_131 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_132 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_133 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_134 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_135 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_136 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_137 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_138 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_139 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_140 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_141 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_142 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_143 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_144 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_145 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_146 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_147 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_148 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_149 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_150 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_151 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_152 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_153 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_154 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_155 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_156 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_157 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_158 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_159 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_160 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_5 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_160 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_159 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_158 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_157 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_156 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_155 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_154 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_153 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_152 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_151 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_150 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_149 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_148 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_147 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_146 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_145 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_144 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_143 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_142 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_141 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_140 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_139 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_138 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_137 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_136 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_135 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_134 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_133 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_132 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_131 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_130 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_129 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_161 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_162 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_163 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_164 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_165 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_166 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_167 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_168 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_169 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_170 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_171 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_172 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_173 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_174 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_175 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_176 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_177 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_178 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_179 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_180 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_181 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_182 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_183 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_184 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_185 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_186 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_187 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_188 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_189 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_190 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_191 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_192 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_6 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_192 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_191 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_190 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_189 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_188 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_187 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_186 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_185 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_184 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_183 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_182 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_181 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_180 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_179 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_178 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_177 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_176 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_175 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_174 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_173 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_172 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_171 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_170 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_169 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_168 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_167 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_166 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_165 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_164 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_163 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_162 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_161 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_3 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_6 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_5 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_193 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_194 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_195 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_196 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_197 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_198 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_199 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_200 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_201 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_202 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_203 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_204 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_205 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_206 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_207 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_208 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_209 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_210 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_211 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_212 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_213 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_214 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_215 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_216 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_217 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_218 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_219 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_220 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_221 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_222 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_223 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_224 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_7 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_224 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_223 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_222 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_221 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_220 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_219 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_218 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_217 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_216 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_215 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_214 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_213 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_212 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_211 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_210 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_209 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_208 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_207 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_206 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_205 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_204 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_203 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_202 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_201 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_200 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_199 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_198 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_197 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_196 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_195 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_194 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_193 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_225 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_226 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_227 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_228 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_229 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_230 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_231 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_232 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_233 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_234 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_235 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_236 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_237 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_238 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_239 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_240 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_241 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_242 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_243 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_244 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_245 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_246 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_247 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_248 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_249 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_250 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_251 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_252 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_253 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_254 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_255 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_256 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_8 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_256 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_255 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_254 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_253 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_252 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_251 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_250 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_249 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_248 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_247 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_246 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_245 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_244 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_243 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_242 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_241 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_240 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_239 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_238 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_237 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_236 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_235 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_234 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_233 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_232 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_231 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_230 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_229 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_228 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_227 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_226 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_225 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_4 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_8 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_7 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_257 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_258 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_259 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_260 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_261 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_262 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_263 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_264 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_265 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_266 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_267 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_268 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_269 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_270 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_271 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_272 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_273 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_274 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_275 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_276 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_277 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_278 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_279 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_280 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_281 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_282 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_283 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_284 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_285 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_286 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_287 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_288 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_9 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_288 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_287 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_286 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_285 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_284 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_283 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_282 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_281 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_280 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_279 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_278 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_277 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_276 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_275 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_274 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_273 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_272 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_271 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_270 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_269 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_268 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_267 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_266 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_265 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_264 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_263 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_262 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_261 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_260 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_259 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_258 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_257 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_289 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_290 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_291 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_292 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_293 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_294 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_295 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_296 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_297 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_298 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_299 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_300 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_301 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_302 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_303 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_304 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_305 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_306 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_307 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_308 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_309 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_310 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_311 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_312 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_313 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_314 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_315 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_316 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_317 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_318 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_319 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_320 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_10 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_320 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_319 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_318 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_317 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_316 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_315 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_314 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_313 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_312 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_311 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_310 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_309 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_308 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_307 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_306 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_305 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_304 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_303 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_302 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_301 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_300 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_299 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_298 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_297 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_296 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_295 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_294 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_293 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_292 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_291 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_290 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_289 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_5 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_10 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_9 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_321 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_322 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_323 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_324 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_325 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_326 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_327 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_328 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_329 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_330 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_331 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_332 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_333 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_334 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_335 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_336 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_337 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_338 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_339 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_340 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_341 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_342 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_343 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_344 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_345 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_346 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_347 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_348 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_349 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_350 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_351 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_352 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_11 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_352 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_351 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_350 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_349 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_348 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_347 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_346 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_345 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_344 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_343 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_342 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_341 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_340 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_339 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_338 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_337 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_336 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_335 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_334 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_333 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_332 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_331 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_330 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_329 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_328 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_327 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_326 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_325 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_324 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_323 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_322 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_321 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_353 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_354 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_355 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_356 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_357 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_358 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_359 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_360 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_361 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_362 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_363 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_364 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_365 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_366 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_367 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_368 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_369 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_370 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_371 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_372 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_373 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_374 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_375 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_376 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_377 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_378 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_379 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_380 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_381 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_382 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_383 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_384 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_12 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_384 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_383 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_382 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_381 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_380 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_379 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_378 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_377 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_376 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_375 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_374 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_373 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_372 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_371 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_370 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_369 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_368 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_367 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_366 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_365 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_364 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_363 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_362 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_361 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_360 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_359 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_358 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_357 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_356 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_355 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_354 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_353 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_6 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_12 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_11 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_385 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_386 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_387 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_388 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_389 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_390 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_391 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_392 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_393 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_394 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_395 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_396 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_397 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_398 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_399 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_400 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_401 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_402 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_403 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_404 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_405 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_406 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_407 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_408 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_409 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_410 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_411 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_412 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_413 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_414 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_415 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_416 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_13 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_416 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_415 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_414 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_413 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_412 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_411 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_410 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_409 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_408 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_407 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_406 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_405 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_404 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_403 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_402 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_401 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_400 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_399 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_398 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_397 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_396 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_395 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_394 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_393 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_392 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_391 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_390 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_389 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_388 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_387 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_386 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_385 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_417 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_418 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_419 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_420 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_421 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_422 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_423 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_424 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_425 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_426 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_427 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_428 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_429 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_430 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_431 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_432 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_433 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_434 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_435 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_436 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_437 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_438 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_439 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_440 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_441 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_442 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_443 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_444 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_445 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_446 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_447 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_448 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_14 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_448 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_447 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_446 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_445 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_444 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_443 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_442 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_441 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_440 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_439 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_438 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_437 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_436 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_435 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_434 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_433 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_432 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_431 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_430 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_429 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_428 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_427 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_426 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_425 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_424 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_423 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_422 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_421 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_420 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_419 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_418 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_417 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_7 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_14 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_13 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_449 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_450 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_451 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_452 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_453 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_454 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_455 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_456 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_457 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_458 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_459 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_460 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_461 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_462 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_463 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_464 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_465 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_466 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_467 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_468 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_469 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_470 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_471 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_472 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_473 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_474 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_475 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_476 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_477 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_478 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_479 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_480 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_15 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_480 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_479 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_478 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_477 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_476 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_475 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_474 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_473 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_472 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_471 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_470 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_469 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_468 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_467 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_466 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_465 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_464 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_463 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_462 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_461 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_460 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_459 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_458 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_457 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_456 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_455 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_454 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_453 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_452 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_451 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_450 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_449 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_481 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_482 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_483 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_484 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_485 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_486 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_487 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_488 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_489 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_490 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_491 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_492 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_493 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_494 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_495 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_496 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_497 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_498 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_499 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_500 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_501 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_502 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_503 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_504 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_505 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_506 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_507 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_508 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_509 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_510 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_511 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_512 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_16 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_512 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_511 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_510 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_509 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_508 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_507 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_506 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_505 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_504 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_503 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_502 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_501 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_500 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_499 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_498 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_497 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_496 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_495 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_494 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_493 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_492 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_491 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_490 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_489 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_488 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_487 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_486 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_485 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_484 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_483 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_482 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_481 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_8 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_16 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_15 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_513 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_514 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_515 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_516 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_517 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_518 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_519 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_520 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_521 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_522 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_523 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_524 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_525 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_526 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_527 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_528 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_529 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_530 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_531 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_532 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_533 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_534 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_535 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_536 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_537 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_538 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_539 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_540 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_541 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_542 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_543 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_544 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_17 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_544 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_543 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_542 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_541 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_540 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_539 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_538 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_537 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_536 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_535 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_534 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_533 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_532 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_531 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_530 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_529 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_528 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_527 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_526 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_525 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_524 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_523 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_522 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_521 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_520 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_519 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_518 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_517 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_516 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_515 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_514 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_513 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_545 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_546 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_547 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_548 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_549 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_550 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_551 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_552 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_553 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_554 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_555 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_556 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_557 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_558 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_559 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_560 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_561 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_562 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_563 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_564 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_565 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_566 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_567 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_568 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_569 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_570 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_571 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_572 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_573 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_574 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_575 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_576 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_18 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_576 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_575 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_574 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_573 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_572 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_571 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_570 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_569 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_568 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_567 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_566 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_565 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_564 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_563 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_562 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_561 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_560 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_559 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_558 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_557 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_556 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_555 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_554 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_553 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_552 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_551 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_550 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_549 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_548 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_547 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_546 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_545 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_9 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_18 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_17 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_577 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_578 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_579 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_580 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_581 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_582 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_583 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_584 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_585 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_586 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_587 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_588 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_589 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_590 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_591 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_592 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_593 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_594 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_595 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_596 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_597 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_598 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_599 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_600 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_601 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_602 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_603 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_604 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_605 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_606 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_607 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_608 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_19 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_608 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_607 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_606 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_605 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_604 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_603 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_602 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_601 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_600 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_599 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_598 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_597 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_596 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_595 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_594 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_593 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_592 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_591 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_590 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_589 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_588 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_587 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_586 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_585 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_584 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_583 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_582 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_581 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_580 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_579 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_578 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_577 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_609 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_610 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_611 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_612 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_613 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_614 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_615 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_616 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_617 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_618 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_619 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_620 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_621 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_622 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_623 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_624 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_625 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_626 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_627 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_628 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_629 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_630 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_631 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_632 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_633 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_634 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_635 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_636 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_637 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_638 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_639 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_640 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_20 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_640 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_639 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_638 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_637 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_636 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_635 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_634 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_633 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_632 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_631 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_630 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_629 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_628 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_627 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_626 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_625 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_624 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_623 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_622 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_621 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_620 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_619 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_618 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_617 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_616 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_615 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_614 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_613 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_612 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_611 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_610 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_609 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_10 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_20 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_19 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_641 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_642 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_643 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_644 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_645 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_646 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_647 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_648 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_649 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_650 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_651 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_652 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_653 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_654 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_655 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_656 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_657 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_658 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_659 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_660 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_661 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_662 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_663 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_664 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_665 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_666 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_667 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_668 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_669 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_670 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_671 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_672 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_21 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_672 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_671 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_670 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_669 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_668 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_667 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_666 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_665 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_664 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_663 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_662 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_661 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_660 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_659 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_658 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_657 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_656 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_655 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_654 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_653 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_652 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_651 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_650 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_649 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_648 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_647 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_646 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_645 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_644 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_643 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_642 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_641 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_673 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_674 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_675 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_676 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_677 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_678 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_679 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_680 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_681 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_682 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_683 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_684 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_685 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_686 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_687 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_688 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_689 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_690 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_691 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_692 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_693 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_694 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_695 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_696 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_697 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_698 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_699 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_700 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_701 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_702 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_703 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_704 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_22 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_704 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_703 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_702 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_701 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_700 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_699 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_698 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_697 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_696 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_695 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_694 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_693 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_692 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_691 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_690 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_689 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_688 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_687 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_686 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_685 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_684 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_683 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_682 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_681 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_680 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_679 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_678 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_677 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_676 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_675 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_674 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_673 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_11 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_22 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_21 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_705 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_706 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_707 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_708 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_709 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_710 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_711 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_712 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_713 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_714 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_715 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_716 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_717 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_718 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_719 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_720 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_721 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_722 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_723 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_724 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_725 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_726 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_727 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_728 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_729 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_730 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_731 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_732 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_733 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_734 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_735 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_736 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_23 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_736 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_735 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_734 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_733 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_732 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_731 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_730 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_729 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_728 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_727 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_726 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_725 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_724 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_723 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_722 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_721 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_720 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_719 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_718 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_717 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_716 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_715 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_714 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_713 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_712 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_711 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_710 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_709 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_708 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_707 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_706 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_705 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_737 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_738 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_739 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_740 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_741 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_742 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_743 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_744 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_745 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_746 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_747 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_748 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_749 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_750 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_751 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_752 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_753 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_754 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_755 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_756 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_757 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_758 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_759 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_760 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_761 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_762 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_763 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_764 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_765 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_766 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_767 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_768 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_24 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_768 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_767 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_766 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_765 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_764 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_763 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_762 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_761 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_760 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_759 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_758 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_757 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_756 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_755 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_754 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_753 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_752 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_751 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_750 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_749 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_748 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_747 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_746 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_745 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_744 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_743 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_742 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_741 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_740 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_739 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_738 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_737 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_12 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_24 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_23 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_769 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_770 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_771 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_772 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_773 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_774 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_775 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_776 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_777 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_778 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_779 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_780 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_781 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_782 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_783 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_784 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_785 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_786 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_787 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_788 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_789 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_790 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_791 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_792 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_793 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_794 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_795 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_796 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_797 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_798 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_799 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_800 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_25 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_800 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_799 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_798 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_797 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_796 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_795 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_794 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_793 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_792 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_791 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_790 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_789 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_788 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_787 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_786 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_785 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_784 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_783 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_782 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_781 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_780 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_779 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_778 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_777 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_776 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_775 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_774 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_773 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_772 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_771 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_770 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_769 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_801 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_802 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_803 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_804 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_805 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_806 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_807 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_808 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_809 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_810 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_811 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_812 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_813 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_814 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_815 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_816 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_817 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_818 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_819 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_820 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_821 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_822 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_823 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_824 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_825 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_826 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_827 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_828 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_829 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_830 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_831 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_832 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_26 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_832 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_831 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_830 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_829 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_828 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_827 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_826 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_825 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_824 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_823 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_822 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_821 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_820 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_819 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_818 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_817 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_816 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_815 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_814 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_813 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_812 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_811 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_810 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_809 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_808 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_807 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_806 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_805 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_804 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_803 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_802 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_801 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_13 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_26 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_25 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_833 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_834 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_835 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_836 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_837 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_838 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_839 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_840 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_841 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_842 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_843 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_844 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_845 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_846 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_847 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_848 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_849 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_850 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_851 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_852 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_853 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_854 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_855 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_856 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_857 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_858 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_859 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_860 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_861 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_862 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_863 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_864 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_27 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_864 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_863 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_862 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_861 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_860 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_859 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_858 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_857 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_856 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_855 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_854 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_853 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_852 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_851 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_850 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_849 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_848 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_847 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_846 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_845 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_844 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_843 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_842 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_841 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_840 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_839 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_838 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_837 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_836 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_835 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_834 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_833 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_865 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_866 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_867 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_868 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_869 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_870 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_871 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_872 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_873 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_874 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_875 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_876 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_877 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_878 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_879 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_880 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_881 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_882 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_883 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_884 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_885 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_886 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_887 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_888 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_889 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_890 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_891 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_892 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_893 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_894 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_895 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_896 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_28 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_896 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_895 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_894 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_893 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_892 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_891 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_890 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_889 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_888 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_887 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_886 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_885 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_884 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_883 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_882 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_881 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_880 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_879 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_878 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_877 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_876 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_875 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_874 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_873 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_872 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_871 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_870 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_869 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_868 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_867 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_866 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_865 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_14 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_28 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_27 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_897 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_898 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_899 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_900 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_901 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_902 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_903 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_904 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_905 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_906 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_907 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_908 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_909 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_910 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_911 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_912 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_913 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_914 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_915 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_916 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_917 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_918 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_919 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_920 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_921 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_922 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_923 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_924 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_925 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_926 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_927 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_928 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_29 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_928 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_927 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_926 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_925 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_924 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_923 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_922 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_921 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_920 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_919 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_918 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_917 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_916 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_915 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_914 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_913 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_912 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_911 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_910 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_909 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_908 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_907 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_906 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_905 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_904 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_903 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_902 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_901 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_900 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_899 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_898 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_897 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_929 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_930 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_931 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_932 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_933 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_934 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_935 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_936 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_937 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_938 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_939 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_940 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_941 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_942 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_943 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_944 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_945 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_946 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_947 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_948 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_949 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_950 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_951 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_952 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_953 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_954 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_955 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_956 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_957 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_958 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_959 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_960 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_30 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_960 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_959 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_958 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_957 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_956 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_955 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_954 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_953 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_952 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_951 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_950 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_949 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_948 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_947 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_946 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_945 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_944 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_943 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_942 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_941 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_940 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_939 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_938 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_937 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_936 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_935 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_934 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_933 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_932 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_931 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_930 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_929 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_15 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_30 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_29 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_961 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_962 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_963 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_964 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_965 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_966 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_967 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_968 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_969 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_970 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_971 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_972 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_973 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_974 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_975 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_976 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_977 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_978 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_979 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_980 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_981 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_982 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_983 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_984 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_985 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_986 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_987 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_988 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_989 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_990 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_991 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_992 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_31 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_992 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_991 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_990 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_989 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_988 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_987 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_986 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_985 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_984 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_983 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_982 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_981 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_980 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_979 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_978 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_977 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_976 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_975 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_974 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_973 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_972 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_971 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_970 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_969 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_968 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_967 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_966 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_965 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_964 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_963 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_962 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_961 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_993 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_994 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_995 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_996 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_997 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_998 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_999 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1000 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1001 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1002 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1003 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1004 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1005 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1006 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1007 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1008 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1009 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1010 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1011 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1012 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1013 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1014 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1015 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1016 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1017 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1018 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1019 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1020 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1021 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1022 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1023 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1024 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_32 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1024 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1023 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1022 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1021 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1020 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1019 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1018 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1017 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1016 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1015 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1014 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1013 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1012 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1011 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1010 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1009 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1008 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1007 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1006 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1005 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1004 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1003 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1002 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1001 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1000 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_999 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_998 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_997 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_996 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_995 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_994 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_993 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_16 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_32 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_31 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1025 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1026 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1027 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1028 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1029 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1030 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1031 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1032 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1033 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1034 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1035 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1036 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1037 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1038 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1039 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1040 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1041 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1042 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1043 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1044 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1045 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1046 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1047 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1048 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1049 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1050 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1051 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1052 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1053 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1054 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1055 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1056 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_33 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1056 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1055 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1054 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1053 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1052 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1051 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1050 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1049 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1048 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1047 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1046 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1045 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1044 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1043 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1042 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1041 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1040 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1039 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1038 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1037 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1036 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1035 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1034 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1033 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1032 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1031 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1030 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1029 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1028 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1027 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1026 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1025 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1057 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1058 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1059 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1060 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1061 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1062 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1063 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1064 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1065 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1066 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1067 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1068 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1069 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1070 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1071 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1072 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1073 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1074 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1075 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1076 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1077 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1078 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1079 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1080 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1081 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1082 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1083 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1084 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1085 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1086 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1087 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1088 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_34 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1088 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1087 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1086 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1085 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1084 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1083 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1082 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1081 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1080 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1079 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1078 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1077 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1076 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1075 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1074 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1073 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1072 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1071 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1070 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1069 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1068 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1067 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1066 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1065 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1064 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1063 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1062 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1061 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1060 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1059 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1058 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1057 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_17 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_34 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_33 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1089 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1090 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1091 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1092 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1093 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1094 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1095 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1096 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1097 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1098 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1099 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1100 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1101 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1102 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1103 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1104 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1105 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1106 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1107 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1108 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1109 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1110 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1111 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1112 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1113 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1114 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1115 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1116 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1117 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1118 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1119 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1120 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_35 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1120 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1119 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1118 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1117 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1116 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1115 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1114 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1113 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1112 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1111 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1110 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1109 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1108 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1107 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1106 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1105 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1104 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1103 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1102 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1101 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1100 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1099 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1098 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1097 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1096 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1095 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1094 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1093 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1092 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1091 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1090 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1089 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1121 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1122 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1123 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1124 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1125 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1126 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1127 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1128 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1129 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1130 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1131 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1132 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1133 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1134 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1135 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1136 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1137 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1138 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1139 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1140 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1141 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1142 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1143 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1144 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1145 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1146 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1147 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1148 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1149 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1150 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1151 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1152 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_36 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1152 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1151 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1150 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1149 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1148 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1147 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1146 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1145 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1144 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1143 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1142 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1141 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1140 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1139 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1138 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1137 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1136 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1135 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1134 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1133 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1132 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1131 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1130 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1129 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1128 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1127 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1126 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1125 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1124 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1123 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1122 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1121 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_18 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_36 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_35 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1153 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1154 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1155 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1156 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1157 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1158 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1159 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1160 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1161 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1162 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1163 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1164 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1165 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1166 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1167 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1168 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1169 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1170 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1171 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1172 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1173 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1174 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1175 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1176 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1177 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1178 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1179 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1180 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1181 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1182 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1183 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1184 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_37 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1184 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1183 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1182 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1181 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1180 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1179 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1178 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1177 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1176 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1175 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1174 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1173 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1172 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1171 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1170 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1169 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1168 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1167 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1166 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1165 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1164 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1163 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1162 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1161 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1160 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1159 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1158 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1157 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1156 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1155 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1154 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1153 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1185 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1186 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1187 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1188 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1189 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1190 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1191 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1192 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1193 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1194 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1195 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1196 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1197 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1198 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1199 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1200 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1201 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1202 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1203 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1204 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1205 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1206 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1207 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1208 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1209 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1210 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1211 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1212 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1213 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1214 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1215 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1216 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_38 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1216 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1215 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1214 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1213 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1212 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1211 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1210 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1209 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1208 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1207 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1206 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1205 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1204 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1203 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1202 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1201 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1200 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1199 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1198 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1197 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1196 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1195 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1194 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1193 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1192 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1191 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1190 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1189 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1188 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1187 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1186 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1185 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_19 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_38 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_37 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1217 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1218 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1219 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1220 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1221 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1222 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1223 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1224 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1225 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1226 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1227 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1228 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1229 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1230 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1231 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1232 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1233 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1234 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1235 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1236 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1237 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1238 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1239 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1240 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1241 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1242 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1243 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1244 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1245 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1246 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1247 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1248 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_39 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1248 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1247 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1246 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1245 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1244 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1243 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1242 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1241 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1240 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1239 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1238 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1237 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1236 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1235 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1234 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1233 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1232 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1231 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1230 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1229 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1228 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1227 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1226 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1225 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1224 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1223 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1222 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1221 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1220 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1219 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1218 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1217 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1249 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1250 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1251 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1252 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1253 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1254 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1255 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1256 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1257 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1258 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1259 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1260 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1261 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1262 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1263 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1264 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1265 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1266 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1267 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1268 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1269 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1270 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1271 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1272 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1273 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1274 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1275 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1276 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1277 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1278 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1279 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1280 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_40 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1280 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1279 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1278 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1277 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1276 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1275 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1274 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1273 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1272 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1271 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1270 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1269 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1268 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1267 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1266 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1265 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1264 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1263 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1262 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1261 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1260 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1259 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1258 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1257 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1256 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1255 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1254 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1253 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1252 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1251 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1250 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1249 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_20 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_40 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_39 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1281 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1282 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1283 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1284 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1285 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1286 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1287 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1288 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1289 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1290 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1291 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1292 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1293 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1294 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1295 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1296 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1297 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1298 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1299 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1300 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1301 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1302 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1303 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1304 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1305 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1306 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1307 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1308 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1309 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1310 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1311 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1312 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_41 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1312 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1311 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1310 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1309 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1308 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1307 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1306 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1305 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1304 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1303 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1302 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1301 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1300 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1299 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1298 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1297 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1296 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1295 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1294 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1293 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1292 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1291 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1290 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1289 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1288 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1287 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1286 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1285 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1284 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1283 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1282 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1281 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1313 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1314 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1315 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1316 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1317 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1318 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1319 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1320 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1321 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1322 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1323 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1324 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1325 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1326 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1327 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1328 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1329 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1330 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1331 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1332 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1333 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1334 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1335 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1336 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1337 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1338 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1339 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1340 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1341 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1342 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1343 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1344 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_42 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1344 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1343 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1342 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1341 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1340 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1339 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1338 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1337 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1336 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1335 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1334 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1333 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1332 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1331 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1330 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1329 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1328 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1327 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1326 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1325 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1324 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1323 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1322 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1321 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1320 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1319 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1318 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1317 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1316 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1315 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1314 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1313 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_21 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_42 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_41 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1345 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1346 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1347 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1348 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1349 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1350 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1351 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1352 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1353 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1354 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1355 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1356 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1357 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1358 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1359 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1360 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1361 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1362 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1363 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1364 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1365 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1366 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1367 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1368 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1369 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1370 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1371 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1372 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1373 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1374 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1375 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1376 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_43 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1376 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1375 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1374 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1373 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1372 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1371 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1370 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1369 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1368 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1367 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1366 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1365 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1364 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1363 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1362 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1361 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1360 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1359 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1358 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1357 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1356 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1355 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1354 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1353 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1352 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1351 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1350 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1349 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1348 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1347 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1346 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1345 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1377 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1378 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1379 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1380 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1381 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1382 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1383 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1384 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1385 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1386 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1387 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1388 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1389 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1390 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1391 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1392 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1393 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1394 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1395 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1396 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1397 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1398 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1399 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1400 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1401 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1402 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1403 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1404 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1405 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1406 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1407 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1408 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_44 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1408 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1407 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1406 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1405 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1404 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1403 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1402 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1401 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1400 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1399 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1398 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1397 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1396 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1395 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1394 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1393 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1392 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1391 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1390 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1389 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1388 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1387 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1386 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1385 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1384 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1383 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1382 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1381 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1380 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1379 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1378 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1377 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_22 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_44 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_43 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1409 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1410 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1411 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1412 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1413 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1414 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1415 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1416 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1417 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1418 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1419 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1420 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1421 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1422 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1423 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1424 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1425 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1426 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1427 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1428 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1429 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1430 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1431 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1432 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1433 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1434 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1435 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1436 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1437 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1438 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1439 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1440 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_45 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1440 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1439 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1438 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1437 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1436 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1435 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1434 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1433 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1432 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1431 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1430 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1429 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1428 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1427 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1426 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1425 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1424 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1423 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1422 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1421 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1420 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1419 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1418 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1417 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1416 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1415 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1414 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1413 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1412 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1411 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1410 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1409 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1441 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1442 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1443 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1444 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1445 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1446 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1447 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1448 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1449 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1450 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1451 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1452 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1453 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1454 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1455 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1456 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1457 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1458 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1459 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1460 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1461 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1462 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1463 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1464 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1465 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1466 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1467 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1468 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1469 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1470 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1471 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1472 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_46 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1472 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1471 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1470 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1469 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1468 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1467 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1466 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1465 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1464 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1463 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1462 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1461 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1460 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1459 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1458 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1457 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1456 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1455 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1454 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1453 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1452 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1451 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1450 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1449 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1448 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1447 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1446 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1445 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1444 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1443 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1442 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1441 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_23 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_46 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_45 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1473 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1474 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1475 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1476 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1477 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1478 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1479 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1480 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1481 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1482 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1483 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1484 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1485 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1486 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1487 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1488 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1489 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1490 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1491 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1492 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1493 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1494 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1495 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1496 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1497 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1498 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1499 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1500 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1501 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1502 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1503 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1504 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_47 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1504 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1503 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1502 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1501 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1500 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1499 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1498 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1497 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1496 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1495 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1494 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1493 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1492 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1491 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1490 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1489 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1488 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1487 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1486 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1485 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1484 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1483 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1482 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1481 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1480 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1479 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1478 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1477 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1476 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1475 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1474 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1473 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1505 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1506 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1507 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1508 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1509 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1510 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1511 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1512 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1513 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1514 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1515 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1516 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1517 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1518 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1519 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1520 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1521 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1522 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1523 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1524 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1525 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1526 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1527 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1528 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1529 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1530 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1531 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1532 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1533 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1534 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1535 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1536 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_48 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1536 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1535 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1534 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1533 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1532 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1531 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1530 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1529 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1528 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1527 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1526 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1525 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1524 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1523 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1522 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1521 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1520 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1519 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1518 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1517 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1516 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1515 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1514 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1513 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1512 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1511 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1510 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1509 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1508 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1507 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1506 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1505 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_24 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_48 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_47 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1537 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1538 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1539 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1540 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1541 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1542 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1543 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1544 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1545 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1546 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1547 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1548 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1549 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1550 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1551 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1552 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1553 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1554 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1555 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1556 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1557 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1558 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1559 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1560 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1561 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1562 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1563 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1564 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1565 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1566 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1567 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1568 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_49 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1568 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1567 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1566 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1565 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1564 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1563 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1562 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1561 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1560 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1559 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1558 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1557 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1556 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1555 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1554 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1553 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1552 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1551 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1550 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1549 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1548 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1547 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1546 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1545 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1544 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1543 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1542 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1541 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1540 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1539 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1538 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1537 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1569 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1570 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1571 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1572 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1573 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1574 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1575 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1576 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1577 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1578 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1579 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1580 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1581 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1582 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1583 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1584 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1585 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1586 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1587 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1588 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1589 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1590 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1591 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1592 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1593 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1594 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1595 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1596 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1597 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1598 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1599 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1600 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_50 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1600 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1599 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1598 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1597 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1596 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1595 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1594 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1593 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1592 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1591 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1590 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1589 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1588 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1587 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1586 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1585 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1584 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1583 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1582 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1581 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1580 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1579 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1578 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1577 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1576 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1575 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1574 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1573 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1572 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1571 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1570 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1569 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_25 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_50 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_49 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1601 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1602 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1603 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1604 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1605 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1606 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1607 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1608 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1609 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1610 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1611 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1612 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1613 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1614 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1615 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1616 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1617 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1618 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1619 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1620 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1621 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1622 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1623 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1624 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1625 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1626 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1627 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1628 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1629 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1630 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1631 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1632 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_51 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1632 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1631 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1630 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1629 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1628 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1627 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1626 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1625 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1624 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1623 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1622 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1621 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1620 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1619 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1618 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1617 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1616 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1615 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1614 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1613 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1612 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1611 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1610 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1609 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1608 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1607 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1606 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1605 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1604 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1603 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1602 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1601 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1633 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1634 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1635 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1636 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1637 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1638 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1639 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1640 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1641 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1642 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1643 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1644 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1645 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1646 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1647 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1648 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1649 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1650 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1651 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1652 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1653 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1654 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1655 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1656 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1657 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1658 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1659 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1660 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1661 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1662 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1663 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1664 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_52 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1664 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1663 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1662 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1661 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1660 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1659 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1658 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1657 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1656 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1655 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1654 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1653 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1652 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1651 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1650 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1649 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1648 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1647 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1646 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1645 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1644 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1643 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1642 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1641 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1640 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1639 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1638 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1637 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1636 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1635 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1634 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1633 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_26 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_52 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_51 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1665 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1666 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1667 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1668 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1669 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1670 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1671 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1672 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1673 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1674 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1675 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1676 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1677 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1678 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1679 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1680 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1681 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1682 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1683 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1684 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1685 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1686 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1687 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1688 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1689 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1690 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1691 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1692 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1693 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1694 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1695 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1696 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_53 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1696 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1695 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1694 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1693 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1692 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1691 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1690 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1689 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1688 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1687 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1686 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1685 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1684 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1683 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1682 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1681 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1680 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1679 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1678 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1677 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1676 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1675 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1674 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1673 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1672 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1671 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1670 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1669 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1668 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1667 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1666 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1665 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1697 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1698 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1699 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1700 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1701 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1702 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1703 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1704 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1705 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1706 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1707 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1708 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1709 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1710 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1711 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1712 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1713 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1714 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1715 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1716 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1717 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1718 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1719 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1720 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1721 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1722 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1723 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1724 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1725 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1726 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1727 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1728 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_54 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1728 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1727 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1726 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1725 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1724 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1723 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1722 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1721 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1720 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1719 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1718 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1717 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1716 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1715 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1714 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1713 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1712 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1711 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1710 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1709 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1708 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1707 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1706 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1705 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1704 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1703 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1702 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1701 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1700 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1699 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1698 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1697 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_27 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_54 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_53 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1729 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1730 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1731 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1732 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1733 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1734 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1735 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1736 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1737 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1738 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1739 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1740 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1741 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1742 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1743 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1744 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1745 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1746 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1747 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1748 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1749 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1750 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1751 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1752 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1753 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1754 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1755 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1756 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1757 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1758 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1759 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1760 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_55 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1760 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1759 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1758 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1757 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1756 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1755 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1754 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1753 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1752 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1751 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1750 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1749 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1748 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1747 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1746 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1745 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1744 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1743 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1742 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1741 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1740 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1739 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1738 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1737 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1736 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1735 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1734 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1733 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1732 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1731 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1730 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1729 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1761 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1762 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1763 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1764 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1765 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1766 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1767 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1768 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1769 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1770 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1771 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1772 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1773 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1774 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1775 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1776 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1777 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1778 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1779 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1780 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1781 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1782 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1783 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1784 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1785 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1786 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1787 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1788 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1789 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1790 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1791 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1792 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_56 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1792 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1791 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1790 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1789 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1788 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1787 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1786 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1785 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1784 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1783 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1782 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1781 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1780 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1779 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1778 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1777 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1776 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1775 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1774 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1773 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1772 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1771 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1770 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1769 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1768 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1767 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1766 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1765 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1764 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1763 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1762 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1761 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_28 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_56 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_55 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1793 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1794 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1795 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1796 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1797 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1798 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1799 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1800 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1801 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1802 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1803 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1804 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1805 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1806 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1807 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1808 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1809 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1810 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1811 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1812 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1813 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1814 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1815 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1816 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1817 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1818 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1819 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1820 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1821 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1822 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1823 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1824 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_57 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1824 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1823 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1822 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1821 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1820 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1819 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1818 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1817 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1816 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1815 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1814 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1813 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1812 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1811 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1810 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1809 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1808 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1807 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1806 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1805 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1804 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1803 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1802 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1801 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1800 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1799 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1798 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1797 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1796 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1795 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1794 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1793 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1825 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1826 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1827 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1828 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1829 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1830 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1831 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1832 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1833 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1834 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1835 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1836 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1837 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1838 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1839 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1840 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1841 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1842 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1843 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1844 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1845 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1846 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1847 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1848 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1849 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1850 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1851 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1852 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1853 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1854 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1855 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1856 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_58 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1856 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1855 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1854 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1853 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1852 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1851 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1850 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1849 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1848 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1847 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1846 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1845 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1844 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1843 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1842 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1841 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1840 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1839 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1838 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1837 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1836 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1835 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1834 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1833 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1832 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1831 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1830 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1829 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1828 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1827 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1826 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1825 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_29 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_58 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_57 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1857 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1858 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1859 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1860 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1861 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1862 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1863 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1864 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1865 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1866 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1867 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1868 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1869 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1870 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1871 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1872 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1873 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1874 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1875 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1876 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1877 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1878 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1879 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1880 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1881 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1882 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1883 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1884 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1885 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1886 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1887 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1888 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_59 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1888 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1887 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1886 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1885 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1884 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1883 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1882 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1881 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1880 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1879 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1878 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1877 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1876 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1875 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1874 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1873 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1872 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1871 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1870 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1869 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1868 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1867 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1866 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1865 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1864 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1863 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1862 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1861 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1860 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1859 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1858 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1857 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1889 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1890 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1891 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1892 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1893 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1894 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1895 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1896 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1897 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1898 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1899 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1900 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1901 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1902 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1903 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1904 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1905 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1906 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1907 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1908 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1909 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1910 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1911 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1912 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1913 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1914 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1915 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1916 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1917 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1918 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1919 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1920 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_60 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1920 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1919 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1918 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1917 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1916 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1915 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1914 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1913 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1912 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1911 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1910 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1909 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1908 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1907 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1906 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1905 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1904 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1903 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1902 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1901 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1900 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1899 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1898 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1897 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1896 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1895 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1894 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1893 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1892 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1891 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1890 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1889 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_30 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_60 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_59 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module FullAdder_1921 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1922 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1923 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1924 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1925 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1926 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1927 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1928 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1929 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1930 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1931 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1932 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1933 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1934 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1935 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1936 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1937 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1938 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1939 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1940 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1941 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1942 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1943 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1944 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1945 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1946 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1947 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1948 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1949 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1950 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1951 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1952 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_61 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1952 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1951 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1950 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1949 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1948 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1947 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1946 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1945 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1944 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1943 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1942 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1941 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1940 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1939 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1938 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1937 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1936 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1935 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1934 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1933 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1932 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1931 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1930 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1929 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1928 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1927 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1926 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1925 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1924 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1923 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1922 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1921 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1953 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1954 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1955 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1956 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1957 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1958 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1959 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1960 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1961 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1962 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1963 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1964 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1965 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1966 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1967 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1968 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1969 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1970 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1971 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1972 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1973 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1974 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1975 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1976 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1977 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1978 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1979 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1980 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1981 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1982 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1983 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1984 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_62 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_1984 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_1983 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_1982 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_1981 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_1980 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_1979 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_1978 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_1977 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_1976 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_1975 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_1974 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_1973 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_1972 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_1971 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_1970 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_1969 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_1968 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_1967 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_1966 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_1965 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_1964 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_1963 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_1962 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_1961 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_1960 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_1959 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_1958 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_1957 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_1956 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_1955 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_1954 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1953 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(
        sum[31]), .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep_31 ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextQ_1 = q[0];
  assign nextA[30] = nextA[31];

  CRAdder_32_62 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_61 sub ( .a(a), .b({n100, n99, n98, n97, n96, n95, n94, n93, n92, 
        n91, n90, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, n79, n78, 
        n77, n76, n75, n74, n73, n72, n71, n70, n69}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U3 ( .A1(n4), .A2(n2), .ZN(n3) );
  NOR2_X4 U4 ( .A1(n68), .A2(q[0]), .ZN(n2) );
  AND2_X2 U5 ( .A1(q[0]), .A2(n68), .ZN(n4) );
  INV_X1 U6 ( .A(n1), .ZN(nextQ[31]) );
  AOI222_X1 U7 ( .A1(sumAM[0]), .A2(n2), .B1(a[0]), .B2(n3), .C1(subAM[0]), 
        .C2(n4), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(nextA[9]) );
  AOI222_X1 U9 ( .A1(sumAM[10]), .A2(n2), .B1(a[10]), .B2(n3), .C1(subAM[10]), 
        .C2(n4), .ZN(n5) );
  INV_X1 U10 ( .A(n6), .ZN(nextA[8]) );
  AOI222_X1 U11 ( .A1(sumAM[9]), .A2(n2), .B1(a[9]), .B2(n3), .C1(subAM[9]), 
        .C2(n4), .ZN(n6) );
  INV_X1 U12 ( .A(n7), .ZN(nextA[7]) );
  AOI222_X1 U13 ( .A1(sumAM[8]), .A2(n2), .B1(a[8]), .B2(n3), .C1(subAM[8]), 
        .C2(n4), .ZN(n7) );
  INV_X1 U14 ( .A(n8), .ZN(nextA[6]) );
  AOI222_X1 U15 ( .A1(sumAM[7]), .A2(n2), .B1(a[7]), .B2(n3), .C1(subAM[7]), 
        .C2(n4), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(nextA[5]) );
  AOI222_X1 U17 ( .A1(sumAM[6]), .A2(n2), .B1(a[6]), .B2(n3), .C1(subAM[6]), 
        .C2(n4), .ZN(n9) );
  INV_X1 U18 ( .A(n10), .ZN(nextA[4]) );
  AOI222_X1 U19 ( .A1(sumAM[5]), .A2(n2), .B1(a[5]), .B2(n3), .C1(subAM[5]), 
        .C2(n4), .ZN(n10) );
  INV_X1 U20 ( .A(n11), .ZN(nextA[3]) );
  AOI222_X1 U21 ( .A1(sumAM[4]), .A2(n2), .B1(a[4]), .B2(n3), .C1(subAM[4]), 
        .C2(n4), .ZN(n11) );
  INV_X1 U22 ( .A(n12), .ZN(nextA[31]) );
  AOI222_X1 U23 ( .A1(sumAM[31]), .A2(n2), .B1(a[31]), .B2(n3), .C1(subAM[31]), 
        .C2(n4), .ZN(n12) );
  INV_X1 U24 ( .A(n13), .ZN(nextA[2]) );
  AOI222_X1 U25 ( .A1(sumAM[3]), .A2(n2), .B1(a[3]), .B2(n3), .C1(subAM[3]), 
        .C2(n4), .ZN(n13) );
  INV_X1 U26 ( .A(n14), .ZN(nextA[29]) );
  AOI222_X1 U27 ( .A1(sumAM[30]), .A2(n2), .B1(a[30]), .B2(n3), .C1(subAM[30]), 
        .C2(n4), .ZN(n14) );
  INV_X1 U28 ( .A(n15), .ZN(nextA[28]) );
  AOI222_X1 U29 ( .A1(sumAM[29]), .A2(n2), .B1(a[29]), .B2(n3), .C1(subAM[29]), 
        .C2(n4), .ZN(n15) );
  INV_X1 U30 ( .A(n16), .ZN(nextA[27]) );
  AOI222_X1 U31 ( .A1(sumAM[28]), .A2(n2), .B1(a[28]), .B2(n3), .C1(subAM[28]), 
        .C2(n4), .ZN(n16) );
  INV_X1 U32 ( .A(n17), .ZN(nextA[26]) );
  AOI222_X1 U33 ( .A1(sumAM[27]), .A2(n2), .B1(a[27]), .B2(n3), .C1(subAM[27]), 
        .C2(n4), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(nextA[25]) );
  AOI222_X1 U35 ( .A1(sumAM[26]), .A2(n2), .B1(a[26]), .B2(n3), .C1(subAM[26]), 
        .C2(n4), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(nextA[24]) );
  AOI222_X1 U37 ( .A1(sumAM[25]), .A2(n2), .B1(a[25]), .B2(n3), .C1(subAM[25]), 
        .C2(n4), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(nextA[23]) );
  AOI222_X1 U39 ( .A1(sumAM[24]), .A2(n2), .B1(a[24]), .B2(n3), .C1(subAM[24]), 
        .C2(n4), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(nextA[22]) );
  AOI222_X1 U41 ( .A1(sumAM[23]), .A2(n2), .B1(a[23]), .B2(n3), .C1(subAM[23]), 
        .C2(n4), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(nextA[21]) );
  AOI222_X1 U43 ( .A1(sumAM[22]), .A2(n2), .B1(a[22]), .B2(n3), .C1(subAM[22]), 
        .C2(n4), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(nextA[20]) );
  AOI222_X1 U45 ( .A1(sumAM[21]), .A2(n2), .B1(a[21]), .B2(n3), .C1(subAM[21]), 
        .C2(n4), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(nextA[1]) );
  AOI222_X1 U47 ( .A1(sumAM[2]), .A2(n2), .B1(a[2]), .B2(n3), .C1(subAM[2]), 
        .C2(n4), .ZN(n24) );
  INV_X1 U48 ( .A(n25), .ZN(nextA[19]) );
  AOI222_X1 U49 ( .A1(sumAM[20]), .A2(n2), .B1(a[20]), .B2(n3), .C1(subAM[20]), 
        .C2(n4), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(nextA[18]) );
  AOI222_X1 U51 ( .A1(sumAM[19]), .A2(n2), .B1(a[19]), .B2(n3), .C1(subAM[19]), 
        .C2(n4), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(nextA[17]) );
  AOI222_X1 U53 ( .A1(sumAM[18]), .A2(n2), .B1(a[18]), .B2(n3), .C1(subAM[18]), 
        .C2(n4), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(nextA[16]) );
  AOI222_X1 U55 ( .A1(sumAM[17]), .A2(n2), .B1(a[17]), .B2(n3), .C1(subAM[17]), 
        .C2(n4), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(nextA[15]) );
  AOI222_X1 U57 ( .A1(sumAM[16]), .A2(n2), .B1(a[16]), .B2(n3), .C1(subAM[16]), 
        .C2(n4), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(nextA[14]) );
  AOI222_X1 U59 ( .A1(sumAM[15]), .A2(n2), .B1(a[15]), .B2(n3), .C1(subAM[15]), 
        .C2(n4), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(nextA[13]) );
  AOI222_X1 U61 ( .A1(sumAM[14]), .A2(n2), .B1(a[14]), .B2(n3), .C1(subAM[14]), 
        .C2(n4), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(nextA[12]) );
  AOI222_X1 U63 ( .A1(sumAM[13]), .A2(n2), .B1(a[13]), .B2(n3), .C1(subAM[13]), 
        .C2(n4), .ZN(n32) );
  INV_X1 U64 ( .A(n65), .ZN(nextA[11]) );
  AOI222_X1 U65 ( .A1(sumAM[12]), .A2(n2), .B1(a[12]), .B2(n3), .C1(subAM[12]), 
        .C2(n4), .ZN(n65) );
  INV_X1 U66 ( .A(n66), .ZN(nextA[10]) );
  AOI222_X1 U67 ( .A1(sumAM[11]), .A2(n2), .B1(a[11]), .B2(n3), .C1(subAM[11]), 
        .C2(n4), .ZN(n66) );
  INV_X1 U68 ( .A(n67), .ZN(nextA[0]) );
  AOI222_X1 U69 ( .A1(sumAM[1]), .A2(n2), .B1(a[1]), .B2(n3), .C1(subAM[1]), 
        .C2(n4), .ZN(n67) );
  INV_X1 U70 ( .A(q_1), .ZN(n68) );
  INV_X1 U71 ( .A(m[0]), .ZN(n69) );
  INV_X1 U72 ( .A(m[1]), .ZN(n70) );
  INV_X1 U73 ( .A(m[2]), .ZN(n71) );
  INV_X1 U74 ( .A(m[3]), .ZN(n72) );
  INV_X1 U75 ( .A(m[4]), .ZN(n73) );
  INV_X1 U76 ( .A(m[5]), .ZN(n74) );
  INV_X1 U77 ( .A(m[6]), .ZN(n75) );
  INV_X1 U78 ( .A(m[7]), .ZN(n76) );
  INV_X1 U79 ( .A(m[8]), .ZN(n77) );
  INV_X1 U80 ( .A(m[9]), .ZN(n78) );
  INV_X1 U81 ( .A(m[10]), .ZN(n79) );
  INV_X1 U82 ( .A(m[11]), .ZN(n80) );
  INV_X1 U83 ( .A(m[12]), .ZN(n81) );
  INV_X1 U84 ( .A(m[13]), .ZN(n82) );
  INV_X1 U85 ( .A(m[14]), .ZN(n83) );
  INV_X1 U86 ( .A(m[15]), .ZN(n84) );
  INV_X1 U87 ( .A(m[16]), .ZN(n85) );
  INV_X1 U88 ( .A(m[17]), .ZN(n86) );
  INV_X1 U89 ( .A(m[18]), .ZN(n87) );
  INV_X1 U90 ( .A(m[19]), .ZN(n88) );
  INV_X1 U91 ( .A(m[20]), .ZN(n89) );
  INV_X1 U92 ( .A(m[21]), .ZN(n90) );
  INV_X1 U93 ( .A(m[22]), .ZN(n91) );
  INV_X1 U94 ( .A(m[23]), .ZN(n92) );
  INV_X1 U95 ( .A(m[24]), .ZN(n93) );
  INV_X1 U96 ( .A(m[25]), .ZN(n94) );
  INV_X1 U97 ( .A(m[26]), .ZN(n95) );
  INV_X1 U98 ( .A(m[27]), .ZN(n96) );
  INV_X1 U99 ( .A(m[28]), .ZN(n97) );
  INV_X1 U100 ( .A(m[29]), .ZN(n98) );
  INV_X1 U101 ( .A(m[30]), .ZN(n99) );
  INV_X1 U102 ( .A(m[31]), .ZN(n100) );
endmodule


module Booth ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;
  wire   nextA_1__31_, nextA_1__30_, nextA_1__29_, nextA_1__28_, nextA_1__27_,
         nextA_1__26_, nextA_1__25_, nextA_1__24_, nextA_1__23_, nextA_1__22_,
         nextA_1__21_, nextA_1__20_, nextA_1__19_, nextA_1__18_, nextA_1__17_,
         nextA_1__16_, nextA_1__15_, nextA_1__14_, nextA_1__13_, nextA_1__12_,
         nextA_1__11_, nextA_1__10_, nextA_1__9_, nextA_1__8_, nextA_1__7_,
         nextA_1__6_, nextA_1__5_, nextA_1__4_, nextA_1__3_, nextA_1__2_,
         nextA_1__1_, nextA_1__0_, nextA_2__31_, nextA_2__30_, nextA_2__29_,
         nextA_2__28_, nextA_2__27_, nextA_2__26_, nextA_2__25_, nextA_2__24_,
         nextA_2__23_, nextA_2__22_, nextA_2__21_, nextA_2__20_, nextA_2__19_,
         nextA_2__18_, nextA_2__17_, nextA_2__16_, nextA_2__15_, nextA_2__14_,
         nextA_2__13_, nextA_2__12_, nextA_2__11_, nextA_2__10_, nextA_2__9_,
         nextA_2__8_, nextA_2__7_, nextA_2__6_, nextA_2__5_, nextA_2__4_,
         nextA_2__3_, nextA_2__2_, nextA_2__1_, nextA_2__0_, nextA_3__31_,
         nextA_3__30_, nextA_3__29_, nextA_3__28_, nextA_3__27_, nextA_3__26_,
         nextA_3__25_, nextA_3__24_, nextA_3__23_, nextA_3__22_, nextA_3__21_,
         nextA_3__20_, nextA_3__19_, nextA_3__18_, nextA_3__17_, nextA_3__16_,
         nextA_3__15_, nextA_3__14_, nextA_3__13_, nextA_3__12_, nextA_3__11_,
         nextA_3__10_, nextA_3__9_, nextA_3__8_, nextA_3__7_, nextA_3__6_,
         nextA_3__5_, nextA_3__4_, nextA_3__3_, nextA_3__2_, nextA_3__1_,
         nextA_3__0_, nextA_4__31_, nextA_4__30_, nextA_4__29_, nextA_4__28_,
         nextA_4__27_, nextA_4__26_, nextA_4__25_, nextA_4__24_, nextA_4__23_,
         nextA_4__22_, nextA_4__21_, nextA_4__20_, nextA_4__19_, nextA_4__18_,
         nextA_4__17_, nextA_4__16_, nextA_4__15_, nextA_4__14_, nextA_4__13_,
         nextA_4__12_, nextA_4__11_, nextA_4__10_, nextA_4__9_, nextA_4__8_,
         nextA_4__7_, nextA_4__6_, nextA_4__5_, nextA_4__4_, nextA_4__3_,
         nextA_4__2_, nextA_4__1_, nextA_4__0_, nextA_5__31_, nextA_5__30_,
         nextA_5__29_, nextA_5__28_, nextA_5__27_, nextA_5__26_, nextA_5__25_,
         nextA_5__24_, nextA_5__23_, nextA_5__22_, nextA_5__21_, nextA_5__20_,
         nextA_5__19_, nextA_5__18_, nextA_5__17_, nextA_5__16_, nextA_5__15_,
         nextA_5__14_, nextA_5__13_, nextA_5__12_, nextA_5__11_, nextA_5__10_,
         nextA_5__9_, nextA_5__8_, nextA_5__7_, nextA_5__6_, nextA_5__5_,
         nextA_5__4_, nextA_5__3_, nextA_5__2_, nextA_5__1_, nextA_5__0_,
         nextA_6__31_, nextA_6__30_, nextA_6__29_, nextA_6__28_, nextA_6__27_,
         nextA_6__26_, nextA_6__25_, nextA_6__24_, nextA_6__23_, nextA_6__22_,
         nextA_6__21_, nextA_6__20_, nextA_6__19_, nextA_6__18_, nextA_6__17_,
         nextA_6__16_, nextA_6__15_, nextA_6__14_, nextA_6__13_, nextA_6__12_,
         nextA_6__11_, nextA_6__10_, nextA_6__9_, nextA_6__8_, nextA_6__7_,
         nextA_6__6_, nextA_6__5_, nextA_6__4_, nextA_6__3_, nextA_6__2_,
         nextA_6__1_, nextA_6__0_, nextA_7__31_, nextA_7__30_, nextA_7__29_,
         nextA_7__28_, nextA_7__27_, nextA_7__26_, nextA_7__25_, nextA_7__24_,
         nextA_7__23_, nextA_7__22_, nextA_7__21_, nextA_7__20_, nextA_7__19_,
         nextA_7__18_, nextA_7__17_, nextA_7__16_, nextA_7__15_, nextA_7__14_,
         nextA_7__13_, nextA_7__12_, nextA_7__11_, nextA_7__10_, nextA_7__9_,
         nextA_7__8_, nextA_7__7_, nextA_7__6_, nextA_7__5_, nextA_7__4_,
         nextA_7__3_, nextA_7__2_, nextA_7__1_, nextA_7__0_, nextA_8__31_,
         nextA_8__30_, nextA_8__29_, nextA_8__28_, nextA_8__27_, nextA_8__26_,
         nextA_8__25_, nextA_8__24_, nextA_8__23_, nextA_8__22_, nextA_8__21_,
         nextA_8__20_, nextA_8__19_, nextA_8__18_, nextA_8__17_, nextA_8__16_,
         nextA_8__15_, nextA_8__14_, nextA_8__13_, nextA_8__12_, nextA_8__11_,
         nextA_8__10_, nextA_8__9_, nextA_8__8_, nextA_8__7_, nextA_8__6_,
         nextA_8__5_, nextA_8__4_, nextA_8__3_, nextA_8__2_, nextA_8__1_,
         nextA_8__0_, nextA_9__31_, nextA_9__30_, nextA_9__29_, nextA_9__28_,
         nextA_9__27_, nextA_9__26_, nextA_9__25_, nextA_9__24_, nextA_9__23_,
         nextA_9__22_, nextA_9__21_, nextA_9__20_, nextA_9__19_, nextA_9__18_,
         nextA_9__17_, nextA_9__16_, nextA_9__15_, nextA_9__14_, nextA_9__13_,
         nextA_9__12_, nextA_9__11_, nextA_9__10_, nextA_9__9_, nextA_9__8_,
         nextA_9__7_, nextA_9__6_, nextA_9__5_, nextA_9__4_, nextA_9__3_,
         nextA_9__2_, nextA_9__1_, nextA_9__0_, nextA_10__31_, nextA_10__30_,
         nextA_10__29_, nextA_10__28_, nextA_10__27_, nextA_10__26_,
         nextA_10__25_, nextA_10__24_, nextA_10__23_, nextA_10__22_,
         nextA_10__21_, nextA_10__20_, nextA_10__19_, nextA_10__18_,
         nextA_10__17_, nextA_10__16_, nextA_10__15_, nextA_10__14_,
         nextA_10__13_, nextA_10__12_, nextA_10__11_, nextA_10__10_,
         nextA_10__9_, nextA_10__8_, nextA_10__7_, nextA_10__6_, nextA_10__5_,
         nextA_10__4_, nextA_10__3_, nextA_10__2_, nextA_10__1_, nextA_10__0_,
         nextA_11__31_, nextA_11__30_, nextA_11__29_, nextA_11__28_,
         nextA_11__27_, nextA_11__26_, nextA_11__25_, nextA_11__24_,
         nextA_11__23_, nextA_11__22_, nextA_11__21_, nextA_11__20_,
         nextA_11__19_, nextA_11__18_, nextA_11__17_, nextA_11__16_,
         nextA_11__15_, nextA_11__14_, nextA_11__13_, nextA_11__12_,
         nextA_11__11_, nextA_11__10_, nextA_11__9_, nextA_11__8_,
         nextA_11__7_, nextA_11__6_, nextA_11__5_, nextA_11__4_, nextA_11__3_,
         nextA_11__2_, nextA_11__1_, nextA_11__0_, nextA_12__31_,
         nextA_12__30_, nextA_12__29_, nextA_12__28_, nextA_12__27_,
         nextA_12__26_, nextA_12__25_, nextA_12__24_, nextA_12__23_,
         nextA_12__22_, nextA_12__21_, nextA_12__20_, nextA_12__19_,
         nextA_12__18_, nextA_12__17_, nextA_12__16_, nextA_12__15_,
         nextA_12__14_, nextA_12__13_, nextA_12__12_, nextA_12__11_,
         nextA_12__10_, nextA_12__9_, nextA_12__8_, nextA_12__7_, nextA_12__6_,
         nextA_12__5_, nextA_12__4_, nextA_12__3_, nextA_12__2_, nextA_12__1_,
         nextA_12__0_, nextA_13__31_, nextA_13__30_, nextA_13__29_,
         nextA_13__28_, nextA_13__27_, nextA_13__26_, nextA_13__25_,
         nextA_13__24_, nextA_13__23_, nextA_13__22_, nextA_13__21_,
         nextA_13__20_, nextA_13__19_, nextA_13__18_, nextA_13__17_,
         nextA_13__16_, nextA_13__15_, nextA_13__14_, nextA_13__13_,
         nextA_13__12_, nextA_13__11_, nextA_13__10_, nextA_13__9_,
         nextA_13__8_, nextA_13__7_, nextA_13__6_, nextA_13__5_, nextA_13__4_,
         nextA_13__3_, nextA_13__2_, nextA_13__1_, nextA_13__0_, nextA_14__31_,
         nextA_14__30_, nextA_14__29_, nextA_14__28_, nextA_14__27_,
         nextA_14__26_, nextA_14__25_, nextA_14__24_, nextA_14__23_,
         nextA_14__22_, nextA_14__21_, nextA_14__20_, nextA_14__19_,
         nextA_14__18_, nextA_14__17_, nextA_14__16_, nextA_14__15_,
         nextA_14__14_, nextA_14__13_, nextA_14__12_, nextA_14__11_,
         nextA_14__10_, nextA_14__9_, nextA_14__8_, nextA_14__7_, nextA_14__6_,
         nextA_14__5_, nextA_14__4_, nextA_14__3_, nextA_14__2_, nextA_14__1_,
         nextA_14__0_, nextA_15__31_, nextA_15__30_, nextA_15__29_,
         nextA_15__28_, nextA_15__27_, nextA_15__26_, nextA_15__25_,
         nextA_15__24_, nextA_15__23_, nextA_15__22_, nextA_15__21_,
         nextA_15__20_, nextA_15__19_, nextA_15__18_, nextA_15__17_,
         nextA_15__16_, nextA_15__15_, nextA_15__14_, nextA_15__13_,
         nextA_15__12_, nextA_15__11_, nextA_15__10_, nextA_15__9_,
         nextA_15__8_, nextA_15__7_, nextA_15__6_, nextA_15__5_, nextA_15__4_,
         nextA_15__3_, nextA_15__2_, nextA_15__1_, nextA_15__0_, nextA_16__31_,
         nextA_16__30_, nextA_16__29_, nextA_16__28_, nextA_16__27_,
         nextA_16__26_, nextA_16__25_, nextA_16__24_, nextA_16__23_,
         nextA_16__22_, nextA_16__21_, nextA_16__20_, nextA_16__19_,
         nextA_16__18_, nextA_16__17_, nextA_16__16_, nextA_16__15_,
         nextA_16__14_, nextA_16__13_, nextA_16__12_, nextA_16__11_,
         nextA_16__10_, nextA_16__9_, nextA_16__8_, nextA_16__7_, nextA_16__6_,
         nextA_16__5_, nextA_16__4_, nextA_16__3_, nextA_16__2_, nextA_16__1_,
         nextA_16__0_, nextA_17__31_, nextA_17__30_, nextA_17__29_,
         nextA_17__28_, nextA_17__27_, nextA_17__26_, nextA_17__25_,
         nextA_17__24_, nextA_17__23_, nextA_17__22_, nextA_17__21_,
         nextA_17__20_, nextA_17__19_, nextA_17__18_, nextA_17__17_,
         nextA_17__16_, nextA_17__15_, nextA_17__14_, nextA_17__13_,
         nextA_17__12_, nextA_17__11_, nextA_17__10_, nextA_17__9_,
         nextA_17__8_, nextA_17__7_, nextA_17__6_, nextA_17__5_, nextA_17__4_,
         nextA_17__3_, nextA_17__2_, nextA_17__1_, nextA_17__0_, nextA_18__31_,
         nextA_18__30_, nextA_18__29_, nextA_18__28_, nextA_18__27_,
         nextA_18__26_, nextA_18__25_, nextA_18__24_, nextA_18__23_,
         nextA_18__22_, nextA_18__21_, nextA_18__20_, nextA_18__19_,
         nextA_18__18_, nextA_18__17_, nextA_18__16_, nextA_18__15_,
         nextA_18__14_, nextA_18__13_, nextA_18__12_, nextA_18__11_,
         nextA_18__10_, nextA_18__9_, nextA_18__8_, nextA_18__7_, nextA_18__6_,
         nextA_18__5_, nextA_18__4_, nextA_18__3_, nextA_18__2_, nextA_18__1_,
         nextA_18__0_, nextA_19__31_, nextA_19__30_, nextA_19__29_,
         nextA_19__28_, nextA_19__27_, nextA_19__26_, nextA_19__25_,
         nextA_19__24_, nextA_19__23_, nextA_19__22_, nextA_19__21_,
         nextA_19__20_, nextA_19__19_, nextA_19__18_, nextA_19__17_,
         nextA_19__16_, nextA_19__15_, nextA_19__14_, nextA_19__13_,
         nextA_19__12_, nextA_19__11_, nextA_19__10_, nextA_19__9_,
         nextA_19__8_, nextA_19__7_, nextA_19__6_, nextA_19__5_, nextA_19__4_,
         nextA_19__3_, nextA_19__2_, nextA_19__1_, nextA_19__0_, nextA_20__31_,
         nextA_20__30_, nextA_20__29_, nextA_20__28_, nextA_20__27_,
         nextA_20__26_, nextA_20__25_, nextA_20__24_, nextA_20__23_,
         nextA_20__22_, nextA_20__21_, nextA_20__20_, nextA_20__19_,
         nextA_20__18_, nextA_20__17_, nextA_20__16_, nextA_20__15_,
         nextA_20__14_, nextA_20__13_, nextA_20__12_, nextA_20__11_,
         nextA_20__10_, nextA_20__9_, nextA_20__8_, nextA_20__7_, nextA_20__6_,
         nextA_20__5_, nextA_20__4_, nextA_20__3_, nextA_20__2_, nextA_20__1_,
         nextA_20__0_, nextA_21__31_, nextA_21__30_, nextA_21__29_,
         nextA_21__28_, nextA_21__27_, nextA_21__26_, nextA_21__25_,
         nextA_21__24_, nextA_21__23_, nextA_21__22_, nextA_21__21_,
         nextA_21__20_, nextA_21__19_, nextA_21__18_, nextA_21__17_,
         nextA_21__16_, nextA_21__15_, nextA_21__14_, nextA_21__13_,
         nextA_21__12_, nextA_21__11_, nextA_21__10_, nextA_21__9_,
         nextA_21__8_, nextA_21__7_, nextA_21__6_, nextA_21__5_, nextA_21__4_,
         nextA_21__3_, nextA_21__2_, nextA_21__1_, nextA_21__0_, nextA_22__31_,
         nextA_22__30_, nextA_22__29_, nextA_22__28_, nextA_22__27_,
         nextA_22__26_, nextA_22__25_, nextA_22__24_, nextA_22__23_,
         nextA_22__22_, nextA_22__21_, nextA_22__20_, nextA_22__19_,
         nextA_22__18_, nextA_22__17_, nextA_22__16_, nextA_22__15_,
         nextA_22__14_, nextA_22__13_, nextA_22__12_, nextA_22__11_,
         nextA_22__10_, nextA_22__9_, nextA_22__8_, nextA_22__7_, nextA_22__6_,
         nextA_22__5_, nextA_22__4_, nextA_22__3_, nextA_22__2_, nextA_22__1_,
         nextA_22__0_, nextA_23__31_, nextA_23__30_, nextA_23__29_,
         nextA_23__28_, nextA_23__27_, nextA_23__26_, nextA_23__25_,
         nextA_23__24_, nextA_23__23_, nextA_23__22_, nextA_23__21_,
         nextA_23__20_, nextA_23__19_, nextA_23__18_, nextA_23__17_,
         nextA_23__16_, nextA_23__15_, nextA_23__14_, nextA_23__13_,
         nextA_23__12_, nextA_23__11_, nextA_23__10_, nextA_23__9_,
         nextA_23__8_, nextA_23__7_, nextA_23__6_, nextA_23__5_, nextA_23__4_,
         nextA_23__3_, nextA_23__2_, nextA_23__1_, nextA_23__0_, nextA_24__31_,
         nextA_24__30_, nextA_24__29_, nextA_24__28_, nextA_24__27_,
         nextA_24__26_, nextA_24__25_, nextA_24__24_, nextA_24__23_,
         nextA_24__22_, nextA_24__21_, nextA_24__20_, nextA_24__19_,
         nextA_24__18_, nextA_24__17_, nextA_24__16_, nextA_24__15_,
         nextA_24__14_, nextA_24__13_, nextA_24__12_, nextA_24__11_,
         nextA_24__10_, nextA_24__9_, nextA_24__8_, nextA_24__7_, nextA_24__6_,
         nextA_24__5_, nextA_24__4_, nextA_24__3_, nextA_24__2_, nextA_24__1_,
         nextA_24__0_, nextA_25__31_, nextA_25__30_, nextA_25__29_,
         nextA_25__28_, nextA_25__27_, nextA_25__26_, nextA_25__25_,
         nextA_25__24_, nextA_25__23_, nextA_25__22_, nextA_25__21_,
         nextA_25__20_, nextA_25__19_, nextA_25__18_, nextA_25__17_,
         nextA_25__16_, nextA_25__15_, nextA_25__14_, nextA_25__13_,
         nextA_25__12_, nextA_25__11_, nextA_25__10_, nextA_25__9_,
         nextA_25__8_, nextA_25__7_, nextA_25__6_, nextA_25__5_, nextA_25__4_,
         nextA_25__3_, nextA_25__2_, nextA_25__1_, nextA_25__0_, nextA_26__31_,
         nextA_26__30_, nextA_26__29_, nextA_26__28_, nextA_26__27_,
         nextA_26__26_, nextA_26__25_, nextA_26__24_, nextA_26__23_,
         nextA_26__22_, nextA_26__21_, nextA_26__20_, nextA_26__19_,
         nextA_26__18_, nextA_26__17_, nextA_26__16_, nextA_26__15_,
         nextA_26__14_, nextA_26__13_, nextA_26__12_, nextA_26__11_,
         nextA_26__10_, nextA_26__9_, nextA_26__8_, nextA_26__7_, nextA_26__6_,
         nextA_26__5_, nextA_26__4_, nextA_26__3_, nextA_26__2_, nextA_26__1_,
         nextA_26__0_, nextA_27__31_, nextA_27__30_, nextA_27__29_,
         nextA_27__28_, nextA_27__27_, nextA_27__26_, nextA_27__25_,
         nextA_27__24_, nextA_27__23_, nextA_27__22_, nextA_27__21_,
         nextA_27__20_, nextA_27__19_, nextA_27__18_, nextA_27__17_,
         nextA_27__16_, nextA_27__15_, nextA_27__14_, nextA_27__13_,
         nextA_27__12_, nextA_27__11_, nextA_27__10_, nextA_27__9_,
         nextA_27__8_, nextA_27__7_, nextA_27__6_, nextA_27__5_, nextA_27__4_,
         nextA_27__3_, nextA_27__2_, nextA_27__1_, nextA_27__0_, nextA_28__31_,
         nextA_28__30_, nextA_28__29_, nextA_28__28_, nextA_28__27_,
         nextA_28__26_, nextA_28__25_, nextA_28__24_, nextA_28__23_,
         nextA_28__22_, nextA_28__21_, nextA_28__20_, nextA_28__19_,
         nextA_28__18_, nextA_28__17_, nextA_28__16_, nextA_28__15_,
         nextA_28__14_, nextA_28__13_, nextA_28__12_, nextA_28__11_,
         nextA_28__10_, nextA_28__9_, nextA_28__8_, nextA_28__7_, nextA_28__6_,
         nextA_28__5_, nextA_28__4_, nextA_28__3_, nextA_28__2_, nextA_28__1_,
         nextA_28__0_, nextA_29__31_, nextA_29__30_, nextA_29__29_,
         nextA_29__28_, nextA_29__27_, nextA_29__26_, nextA_29__25_,
         nextA_29__24_, nextA_29__23_, nextA_29__22_, nextA_29__21_,
         nextA_29__20_, nextA_29__19_, nextA_29__18_, nextA_29__17_,
         nextA_29__16_, nextA_29__15_, nextA_29__14_, nextA_29__13_,
         nextA_29__12_, nextA_29__11_, nextA_29__10_, nextA_29__9_,
         nextA_29__8_, nextA_29__7_, nextA_29__6_, nextA_29__5_, nextA_29__4_,
         nextA_29__3_, nextA_29__2_, nextA_29__1_, nextA_29__0_, nextA_30__31_,
         nextA_30__30_, nextA_30__29_, nextA_30__28_, nextA_30__27_,
         nextA_30__26_, nextA_30__25_, nextA_30__24_, nextA_30__23_,
         nextA_30__22_, nextA_30__21_, nextA_30__20_, nextA_30__19_,
         nextA_30__18_, nextA_30__17_, nextA_30__16_, nextA_30__15_,
         nextA_30__14_, nextA_30__13_, nextA_30__12_, nextA_30__11_,
         nextA_30__10_, nextA_30__9_, nextA_30__8_, nextA_30__7_, nextA_30__6_,
         nextA_30__5_, nextA_30__4_, nextA_30__3_, nextA_30__2_, nextA_30__1_,
         nextA_30__0_, nextA_31__31_, nextA_31__30_, nextA_31__29_,
         nextA_31__28_, nextA_31__27_, nextA_31__26_, nextA_31__25_,
         nextA_31__24_, nextA_31__23_, nextA_31__22_, nextA_31__21_,
         nextA_31__20_, nextA_31__19_, nextA_31__18_, nextA_31__17_,
         nextA_31__16_, nextA_31__15_, nextA_31__14_, nextA_31__13_,
         nextA_31__12_, nextA_31__11_, nextA_31__10_, nextA_31__9_,
         nextA_31__8_, nextA_31__7_, nextA_31__6_, nextA_31__5_, nextA_31__4_,
         nextA_31__3_, nextA_31__2_, nextA_31__1_, nextA_31__0_, nextQ_1__31_,
         nextQ_1__30_, nextQ_1__29_, nextQ_1__28_, nextQ_1__27_, nextQ_1__26_,
         nextQ_1__25_, nextQ_1__24_, nextQ_1__23_, nextQ_1__22_, nextQ_1__21_,
         nextQ_1__20_, nextQ_1__19_, nextQ_1__18_, nextQ_1__17_, nextQ_1__16_,
         nextQ_1__15_, nextQ_1__14_, nextQ_1__13_, nextQ_1__12_, nextQ_1__11_,
         nextQ_1__10_, nextQ_1__9_, nextQ_1__8_, nextQ_1__7_, nextQ_1__6_,
         nextQ_1__5_, nextQ_1__4_, nextQ_1__3_, nextQ_1__2_, nextQ_1__1_,
         nextQ_1__0_, nextQ_2__31_, nextQ_2__30_, nextQ_2__29_, nextQ_2__28_,
         nextQ_2__27_, nextQ_2__26_, nextQ_2__25_, nextQ_2__24_, nextQ_2__23_,
         nextQ_2__22_, nextQ_2__21_, nextQ_2__20_, nextQ_2__19_, nextQ_2__18_,
         nextQ_2__17_, nextQ_2__16_, nextQ_2__15_, nextQ_2__14_, nextQ_2__13_,
         nextQ_2__12_, nextQ_2__11_, nextQ_2__10_, nextQ_2__9_, nextQ_2__8_,
         nextQ_2__7_, nextQ_2__6_, nextQ_2__5_, nextQ_2__4_, nextQ_2__3_,
         nextQ_2__2_, nextQ_2__1_, nextQ_2__0_, nextQ_3__31_, nextQ_3__30_,
         nextQ_3__29_, nextQ_3__28_, nextQ_3__27_, nextQ_3__26_, nextQ_3__25_,
         nextQ_3__24_, nextQ_3__23_, nextQ_3__22_, nextQ_3__21_, nextQ_3__20_,
         nextQ_3__19_, nextQ_3__18_, nextQ_3__17_, nextQ_3__16_, nextQ_3__15_,
         nextQ_3__14_, nextQ_3__13_, nextQ_3__12_, nextQ_3__11_, nextQ_3__10_,
         nextQ_3__9_, nextQ_3__8_, nextQ_3__7_, nextQ_3__6_, nextQ_3__5_,
         nextQ_3__4_, nextQ_3__3_, nextQ_3__2_, nextQ_3__1_, nextQ_3__0_,
         nextQ_4__31_, nextQ_4__30_, nextQ_4__29_, nextQ_4__28_, nextQ_4__27_,
         nextQ_4__26_, nextQ_4__25_, nextQ_4__24_, nextQ_4__23_, nextQ_4__22_,
         nextQ_4__21_, nextQ_4__20_, nextQ_4__19_, nextQ_4__18_, nextQ_4__17_,
         nextQ_4__16_, nextQ_4__15_, nextQ_4__14_, nextQ_4__13_, nextQ_4__12_,
         nextQ_4__11_, nextQ_4__10_, nextQ_4__9_, nextQ_4__8_, nextQ_4__7_,
         nextQ_4__6_, nextQ_4__5_, nextQ_4__4_, nextQ_4__3_, nextQ_4__2_,
         nextQ_4__1_, nextQ_4__0_, nextQ_5__31_, nextQ_5__30_, nextQ_5__29_,
         nextQ_5__28_, nextQ_5__27_, nextQ_5__26_, nextQ_5__25_, nextQ_5__24_,
         nextQ_5__23_, nextQ_5__22_, nextQ_5__21_, nextQ_5__20_, nextQ_5__19_,
         nextQ_5__18_, nextQ_5__17_, nextQ_5__16_, nextQ_5__15_, nextQ_5__14_,
         nextQ_5__13_, nextQ_5__12_, nextQ_5__11_, nextQ_5__10_, nextQ_5__9_,
         nextQ_5__8_, nextQ_5__7_, nextQ_5__6_, nextQ_5__5_, nextQ_5__4_,
         nextQ_5__3_, nextQ_5__2_, nextQ_5__1_, nextQ_5__0_, nextQ_6__31_,
         nextQ_6__30_, nextQ_6__29_, nextQ_6__28_, nextQ_6__27_, nextQ_6__26_,
         nextQ_6__25_, nextQ_6__24_, nextQ_6__23_, nextQ_6__22_, nextQ_6__21_,
         nextQ_6__20_, nextQ_6__19_, nextQ_6__18_, nextQ_6__17_, nextQ_6__16_,
         nextQ_6__15_, nextQ_6__14_, nextQ_6__13_, nextQ_6__12_, nextQ_6__11_,
         nextQ_6__10_, nextQ_6__9_, nextQ_6__8_, nextQ_6__7_, nextQ_6__6_,
         nextQ_6__5_, nextQ_6__4_, nextQ_6__3_, nextQ_6__2_, nextQ_6__1_,
         nextQ_6__0_, nextQ_7__31_, nextQ_7__30_, nextQ_7__29_, nextQ_7__28_,
         nextQ_7__27_, nextQ_7__26_, nextQ_7__25_, nextQ_7__24_, nextQ_7__23_,
         nextQ_7__22_, nextQ_7__21_, nextQ_7__20_, nextQ_7__19_, nextQ_7__18_,
         nextQ_7__17_, nextQ_7__16_, nextQ_7__15_, nextQ_7__14_, nextQ_7__13_,
         nextQ_7__12_, nextQ_7__11_, nextQ_7__10_, nextQ_7__9_, nextQ_7__8_,
         nextQ_7__7_, nextQ_7__6_, nextQ_7__5_, nextQ_7__4_, nextQ_7__3_,
         nextQ_7__2_, nextQ_7__1_, nextQ_7__0_, nextQ_8__31_, nextQ_8__30_,
         nextQ_8__29_, nextQ_8__28_, nextQ_8__27_, nextQ_8__26_, nextQ_8__25_,
         nextQ_8__24_, nextQ_8__23_, nextQ_8__22_, nextQ_8__21_, nextQ_8__20_,
         nextQ_8__19_, nextQ_8__18_, nextQ_8__17_, nextQ_8__16_, nextQ_8__15_,
         nextQ_8__14_, nextQ_8__13_, nextQ_8__12_, nextQ_8__11_, nextQ_8__10_,
         nextQ_8__9_, nextQ_8__8_, nextQ_8__7_, nextQ_8__6_, nextQ_8__5_,
         nextQ_8__4_, nextQ_8__3_, nextQ_8__2_, nextQ_8__1_, nextQ_8__0_,
         nextQ_9__31_, nextQ_9__30_, nextQ_9__29_, nextQ_9__28_, nextQ_9__27_,
         nextQ_9__26_, nextQ_9__25_, nextQ_9__24_, nextQ_9__23_, nextQ_9__22_,
         nextQ_9__21_, nextQ_9__20_, nextQ_9__19_, nextQ_9__18_, nextQ_9__17_,
         nextQ_9__16_, nextQ_9__15_, nextQ_9__14_, nextQ_9__13_, nextQ_9__12_,
         nextQ_9__11_, nextQ_9__10_, nextQ_9__9_, nextQ_9__8_, nextQ_9__7_,
         nextQ_9__6_, nextQ_9__5_, nextQ_9__4_, nextQ_9__3_, nextQ_9__2_,
         nextQ_9__1_, nextQ_9__0_, nextQ_10__31_, nextQ_10__30_, nextQ_10__29_,
         nextQ_10__28_, nextQ_10__27_, nextQ_10__26_, nextQ_10__25_,
         nextQ_10__24_, nextQ_10__23_, nextQ_10__22_, nextQ_10__21_,
         nextQ_10__20_, nextQ_10__19_, nextQ_10__18_, nextQ_10__17_,
         nextQ_10__16_, nextQ_10__15_, nextQ_10__14_, nextQ_10__13_,
         nextQ_10__12_, nextQ_10__11_, nextQ_10__10_, nextQ_10__9_,
         nextQ_10__8_, nextQ_10__7_, nextQ_10__6_, nextQ_10__5_, nextQ_10__4_,
         nextQ_10__3_, nextQ_10__2_, nextQ_10__1_, nextQ_10__0_, nextQ_11__31_,
         nextQ_11__30_, nextQ_11__29_, nextQ_11__28_, nextQ_11__27_,
         nextQ_11__26_, nextQ_11__25_, nextQ_11__24_, nextQ_11__23_,
         nextQ_11__22_, nextQ_11__21_, nextQ_11__20_, nextQ_11__19_,
         nextQ_11__18_, nextQ_11__17_, nextQ_11__16_, nextQ_11__15_,
         nextQ_11__14_, nextQ_11__13_, nextQ_11__12_, nextQ_11__11_,
         nextQ_11__10_, nextQ_11__9_, nextQ_11__8_, nextQ_11__7_, nextQ_11__6_,
         nextQ_11__5_, nextQ_11__4_, nextQ_11__3_, nextQ_11__2_, nextQ_11__1_,
         nextQ_11__0_, nextQ_12__31_, nextQ_12__30_, nextQ_12__29_,
         nextQ_12__28_, nextQ_12__27_, nextQ_12__26_, nextQ_12__25_,
         nextQ_12__24_, nextQ_12__23_, nextQ_12__22_, nextQ_12__21_,
         nextQ_12__20_, nextQ_12__19_, nextQ_12__18_, nextQ_12__17_,
         nextQ_12__16_, nextQ_12__15_, nextQ_12__14_, nextQ_12__13_,
         nextQ_12__12_, nextQ_12__11_, nextQ_12__10_, nextQ_12__9_,
         nextQ_12__8_, nextQ_12__7_, nextQ_12__6_, nextQ_12__5_, nextQ_12__4_,
         nextQ_12__3_, nextQ_12__2_, nextQ_12__1_, nextQ_12__0_, nextQ_13__31_,
         nextQ_13__30_, nextQ_13__29_, nextQ_13__28_, nextQ_13__27_,
         nextQ_13__26_, nextQ_13__25_, nextQ_13__24_, nextQ_13__23_,
         nextQ_13__22_, nextQ_13__21_, nextQ_13__20_, nextQ_13__19_,
         nextQ_13__18_, nextQ_13__17_, nextQ_13__16_, nextQ_13__15_,
         nextQ_13__14_, nextQ_13__13_, nextQ_13__12_, nextQ_13__11_,
         nextQ_13__10_, nextQ_13__9_, nextQ_13__8_, nextQ_13__7_, nextQ_13__6_,
         nextQ_13__5_, nextQ_13__4_, nextQ_13__3_, nextQ_13__2_, nextQ_13__1_,
         nextQ_13__0_, nextQ_14__31_, nextQ_14__30_, nextQ_14__29_,
         nextQ_14__28_, nextQ_14__27_, nextQ_14__26_, nextQ_14__25_,
         nextQ_14__24_, nextQ_14__23_, nextQ_14__22_, nextQ_14__21_,
         nextQ_14__20_, nextQ_14__19_, nextQ_14__18_, nextQ_14__17_,
         nextQ_14__16_, nextQ_14__15_, nextQ_14__14_, nextQ_14__13_,
         nextQ_14__12_, nextQ_14__11_, nextQ_14__10_, nextQ_14__9_,
         nextQ_14__8_, nextQ_14__7_, nextQ_14__6_, nextQ_14__5_, nextQ_14__4_,
         nextQ_14__3_, nextQ_14__2_, nextQ_14__1_, nextQ_14__0_, nextQ_15__31_,
         nextQ_15__30_, nextQ_15__29_, nextQ_15__28_, nextQ_15__27_,
         nextQ_15__26_, nextQ_15__25_, nextQ_15__24_, nextQ_15__23_,
         nextQ_15__22_, nextQ_15__21_, nextQ_15__20_, nextQ_15__19_,
         nextQ_15__18_, nextQ_15__17_, nextQ_15__16_, nextQ_15__15_,
         nextQ_15__14_, nextQ_15__13_, nextQ_15__12_, nextQ_15__11_,
         nextQ_15__10_, nextQ_15__9_, nextQ_15__8_, nextQ_15__7_, nextQ_15__6_,
         nextQ_15__5_, nextQ_15__4_, nextQ_15__3_, nextQ_15__2_, nextQ_15__1_,
         nextQ_15__0_, nextQ_16__31_, nextQ_16__30_, nextQ_16__29_,
         nextQ_16__28_, nextQ_16__27_, nextQ_16__26_, nextQ_16__25_,
         nextQ_16__24_, nextQ_16__23_, nextQ_16__22_, nextQ_16__21_,
         nextQ_16__20_, nextQ_16__19_, nextQ_16__18_, nextQ_16__17_,
         nextQ_16__16_, nextQ_16__15_, nextQ_16__14_, nextQ_16__13_,
         nextQ_16__12_, nextQ_16__11_, nextQ_16__10_, nextQ_16__9_,
         nextQ_16__8_, nextQ_16__7_, nextQ_16__6_, nextQ_16__5_, nextQ_16__4_,
         nextQ_16__3_, nextQ_16__2_, nextQ_16__1_, nextQ_16__0_, nextQ_17__31_,
         nextQ_17__30_, nextQ_17__29_, nextQ_17__28_, nextQ_17__27_,
         nextQ_17__26_, nextQ_17__25_, nextQ_17__24_, nextQ_17__23_,
         nextQ_17__22_, nextQ_17__21_, nextQ_17__20_, nextQ_17__19_,
         nextQ_17__18_, nextQ_17__17_, nextQ_17__16_, nextQ_17__15_,
         nextQ_17__14_, nextQ_17__13_, nextQ_17__12_, nextQ_17__11_,
         nextQ_17__10_, nextQ_17__9_, nextQ_17__8_, nextQ_17__7_, nextQ_17__6_,
         nextQ_17__5_, nextQ_17__4_, nextQ_17__3_, nextQ_17__2_, nextQ_17__1_,
         nextQ_17__0_, nextQ_18__31_, nextQ_18__30_, nextQ_18__29_,
         nextQ_18__28_, nextQ_18__27_, nextQ_18__26_, nextQ_18__25_,
         nextQ_18__24_, nextQ_18__23_, nextQ_18__22_, nextQ_18__21_,
         nextQ_18__20_, nextQ_18__19_, nextQ_18__18_, nextQ_18__17_,
         nextQ_18__16_, nextQ_18__15_, nextQ_18__14_, nextQ_18__13_,
         nextQ_18__12_, nextQ_18__11_, nextQ_18__10_, nextQ_18__9_,
         nextQ_18__8_, nextQ_18__7_, nextQ_18__6_, nextQ_18__5_, nextQ_18__4_,
         nextQ_18__3_, nextQ_18__2_, nextQ_18__1_, nextQ_18__0_, nextQ_19__31_,
         nextQ_19__30_, nextQ_19__29_, nextQ_19__28_, nextQ_19__27_,
         nextQ_19__26_, nextQ_19__25_, nextQ_19__24_, nextQ_19__23_,
         nextQ_19__22_, nextQ_19__21_, nextQ_19__20_, nextQ_19__19_,
         nextQ_19__18_, nextQ_19__17_, nextQ_19__16_, nextQ_19__15_,
         nextQ_19__14_, nextQ_19__13_, nextQ_19__12_, nextQ_19__11_,
         nextQ_19__10_, nextQ_19__9_, nextQ_19__8_, nextQ_19__7_, nextQ_19__6_,
         nextQ_19__5_, nextQ_19__4_, nextQ_19__3_, nextQ_19__2_, nextQ_19__1_,
         nextQ_19__0_, nextQ_20__31_, nextQ_20__30_, nextQ_20__29_,
         nextQ_20__28_, nextQ_20__27_, nextQ_20__26_, nextQ_20__25_,
         nextQ_20__24_, nextQ_20__23_, nextQ_20__22_, nextQ_20__21_,
         nextQ_20__20_, nextQ_20__19_, nextQ_20__18_, nextQ_20__17_,
         nextQ_20__16_, nextQ_20__15_, nextQ_20__14_, nextQ_20__13_,
         nextQ_20__12_, nextQ_20__11_, nextQ_20__10_, nextQ_20__9_,
         nextQ_20__8_, nextQ_20__7_, nextQ_20__6_, nextQ_20__5_, nextQ_20__4_,
         nextQ_20__3_, nextQ_20__2_, nextQ_20__1_, nextQ_20__0_, nextQ_21__31_,
         nextQ_21__30_, nextQ_21__29_, nextQ_21__28_, nextQ_21__27_,
         nextQ_21__26_, nextQ_21__25_, nextQ_21__24_, nextQ_21__23_,
         nextQ_21__22_, nextQ_21__21_, nextQ_21__20_, nextQ_21__19_,
         nextQ_21__18_, nextQ_21__17_, nextQ_21__16_, nextQ_21__15_,
         nextQ_21__14_, nextQ_21__13_, nextQ_21__12_, nextQ_21__11_,
         nextQ_21__10_, nextQ_21__9_, nextQ_21__8_, nextQ_21__7_, nextQ_21__6_,
         nextQ_21__5_, nextQ_21__4_, nextQ_21__3_, nextQ_21__2_, nextQ_21__1_,
         nextQ_21__0_, nextQ_22__31_, nextQ_22__30_, nextQ_22__29_,
         nextQ_22__28_, nextQ_22__27_, nextQ_22__26_, nextQ_22__25_,
         nextQ_22__24_, nextQ_22__23_, nextQ_22__22_, nextQ_22__21_,
         nextQ_22__20_, nextQ_22__19_, nextQ_22__18_, nextQ_22__17_,
         nextQ_22__16_, nextQ_22__15_, nextQ_22__14_, nextQ_22__13_,
         nextQ_22__12_, nextQ_22__11_, nextQ_22__10_, nextQ_22__9_,
         nextQ_22__8_, nextQ_22__7_, nextQ_22__6_, nextQ_22__5_, nextQ_22__4_,
         nextQ_22__3_, nextQ_22__2_, nextQ_22__1_, nextQ_22__0_, nextQ_23__31_,
         nextQ_23__30_, nextQ_23__29_, nextQ_23__28_, nextQ_23__27_,
         nextQ_23__26_, nextQ_23__25_, nextQ_23__24_, nextQ_23__23_,
         nextQ_23__22_, nextQ_23__21_, nextQ_23__20_, nextQ_23__19_,
         nextQ_23__18_, nextQ_23__17_, nextQ_23__16_, nextQ_23__15_,
         nextQ_23__14_, nextQ_23__13_, nextQ_23__12_, nextQ_23__11_,
         nextQ_23__10_, nextQ_23__9_, nextQ_23__8_, nextQ_23__7_, nextQ_23__6_,
         nextQ_23__5_, nextQ_23__4_, nextQ_23__3_, nextQ_23__2_, nextQ_23__1_,
         nextQ_23__0_, nextQ_24__31_, nextQ_24__30_, nextQ_24__29_,
         nextQ_24__28_, nextQ_24__27_, nextQ_24__26_, nextQ_24__25_,
         nextQ_24__24_, nextQ_24__23_, nextQ_24__22_, nextQ_24__21_,
         nextQ_24__20_, nextQ_24__19_, nextQ_24__18_, nextQ_24__17_,
         nextQ_24__16_, nextQ_24__15_, nextQ_24__14_, nextQ_24__13_,
         nextQ_24__12_, nextQ_24__11_, nextQ_24__10_, nextQ_24__9_,
         nextQ_24__8_, nextQ_24__7_, nextQ_24__6_, nextQ_24__5_, nextQ_24__4_,
         nextQ_24__3_, nextQ_24__2_, nextQ_24__1_, nextQ_24__0_, nextQ_25__31_,
         nextQ_25__30_, nextQ_25__29_, nextQ_25__28_, nextQ_25__27_,
         nextQ_25__26_, nextQ_25__25_, nextQ_25__24_, nextQ_25__23_,
         nextQ_25__22_, nextQ_25__21_, nextQ_25__20_, nextQ_25__19_,
         nextQ_25__18_, nextQ_25__17_, nextQ_25__16_, nextQ_25__15_,
         nextQ_25__14_, nextQ_25__13_, nextQ_25__12_, nextQ_25__11_,
         nextQ_25__10_, nextQ_25__9_, nextQ_25__8_, nextQ_25__7_, nextQ_25__6_,
         nextQ_25__5_, nextQ_25__4_, nextQ_25__3_, nextQ_25__2_, nextQ_25__1_,
         nextQ_25__0_, nextQ_26__31_, nextQ_26__30_, nextQ_26__29_,
         nextQ_26__28_, nextQ_26__27_, nextQ_26__26_, nextQ_26__25_,
         nextQ_26__24_, nextQ_26__23_, nextQ_26__22_, nextQ_26__21_,
         nextQ_26__20_, nextQ_26__19_, nextQ_26__18_, nextQ_26__17_,
         nextQ_26__16_, nextQ_26__15_, nextQ_26__14_, nextQ_26__13_,
         nextQ_26__12_, nextQ_26__11_, nextQ_26__10_, nextQ_26__9_,
         nextQ_26__8_, nextQ_26__7_, nextQ_26__6_, nextQ_26__5_, nextQ_26__4_,
         nextQ_26__3_, nextQ_26__2_, nextQ_26__1_, nextQ_26__0_, nextQ_27__31_,
         nextQ_27__30_, nextQ_27__29_, nextQ_27__28_, nextQ_27__27_,
         nextQ_27__26_, nextQ_27__25_, nextQ_27__24_, nextQ_27__23_,
         nextQ_27__22_, nextQ_27__21_, nextQ_27__20_, nextQ_27__19_,
         nextQ_27__18_, nextQ_27__17_, nextQ_27__16_, nextQ_27__15_,
         nextQ_27__14_, nextQ_27__13_, nextQ_27__12_, nextQ_27__11_,
         nextQ_27__10_, nextQ_27__9_, nextQ_27__8_, nextQ_27__7_, nextQ_27__6_,
         nextQ_27__5_, nextQ_27__4_, nextQ_27__3_, nextQ_27__2_, nextQ_27__1_,
         nextQ_27__0_, nextQ_28__31_, nextQ_28__30_, nextQ_28__29_,
         nextQ_28__28_, nextQ_28__27_, nextQ_28__26_, nextQ_28__25_,
         nextQ_28__24_, nextQ_28__23_, nextQ_28__22_, nextQ_28__21_,
         nextQ_28__20_, nextQ_28__19_, nextQ_28__18_, nextQ_28__17_,
         nextQ_28__16_, nextQ_28__15_, nextQ_28__14_, nextQ_28__13_,
         nextQ_28__12_, nextQ_28__11_, nextQ_28__10_, nextQ_28__9_,
         nextQ_28__8_, nextQ_28__7_, nextQ_28__6_, nextQ_28__5_, nextQ_28__4_,
         nextQ_28__3_, nextQ_28__2_, nextQ_28__1_, nextQ_28__0_, nextQ_29__31_,
         nextQ_29__30_, nextQ_29__29_, nextQ_29__28_, nextQ_29__27_,
         nextQ_29__26_, nextQ_29__25_, nextQ_29__24_, nextQ_29__23_,
         nextQ_29__22_, nextQ_29__21_, nextQ_29__20_, nextQ_29__19_,
         nextQ_29__18_, nextQ_29__17_, nextQ_29__16_, nextQ_29__15_,
         nextQ_29__14_, nextQ_29__13_, nextQ_29__12_, nextQ_29__11_,
         nextQ_29__10_, nextQ_29__9_, nextQ_29__8_, nextQ_29__7_, nextQ_29__6_,
         nextQ_29__5_, nextQ_29__4_, nextQ_29__3_, nextQ_29__2_, nextQ_29__1_,
         nextQ_29__0_, nextQ_30__31_, nextQ_30__30_, nextQ_30__29_,
         nextQ_30__28_, nextQ_30__27_, nextQ_30__26_, nextQ_30__25_,
         nextQ_30__24_, nextQ_30__23_, nextQ_30__22_, nextQ_30__21_,
         nextQ_30__20_, nextQ_30__19_, nextQ_30__18_, nextQ_30__17_,
         nextQ_30__16_, nextQ_30__15_, nextQ_30__14_, nextQ_30__13_,
         nextQ_30__12_, nextQ_30__11_, nextQ_30__10_, nextQ_30__9_,
         nextQ_30__8_, nextQ_30__7_, nextQ_30__6_, nextQ_30__5_, nextQ_30__4_,
         nextQ_30__3_, nextQ_30__2_, nextQ_30__1_, nextQ_30__0_, nextQ_31__31_,
         nextQ_31__30_, nextQ_31__29_, nextQ_31__28_, nextQ_31__27_,
         nextQ_31__26_, nextQ_31__25_, nextQ_31__24_, nextQ_31__23_,
         nextQ_31__22_, nextQ_31__21_, nextQ_31__20_, nextQ_31__19_,
         nextQ_31__18_, nextQ_31__17_, nextQ_31__16_, nextQ_31__15_,
         nextQ_31__14_, nextQ_31__13_, nextQ_31__12_, nextQ_31__11_,
         nextQ_31__10_, nextQ_31__9_, nextQ_31__8_, nextQ_31__7_, nextQ_31__6_,
         nextQ_31__5_, nextQ_31__4_, nextQ_31__3_, nextQ_31__2_, nextQ_31__1_,
         nextQ_31__0_;
  wire   [31:1] q_1;

  BoothStep_0 booth_instances_0__stepX ( .a({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .q(b), .m(a), .q_1(1'b0), .nextA({nextA_1__31_, 
        nextA_1__30_, nextA_1__29_, nextA_1__28_, nextA_1__27_, nextA_1__26_, 
        nextA_1__25_, nextA_1__24_, nextA_1__23_, nextA_1__22_, nextA_1__21_, 
        nextA_1__20_, nextA_1__19_, nextA_1__18_, nextA_1__17_, nextA_1__16_, 
        nextA_1__15_, nextA_1__14_, nextA_1__13_, nextA_1__12_, nextA_1__11_, 
        nextA_1__10_, nextA_1__9_, nextA_1__8_, nextA_1__7_, nextA_1__6_, 
        nextA_1__5_, nextA_1__4_, nextA_1__3_, nextA_1__2_, nextA_1__1_, 
        nextA_1__0_}), .nextQ({nextQ_1__31_, nextQ_1__30_, nextQ_1__29_, 
        nextQ_1__28_, nextQ_1__27_, nextQ_1__26_, nextQ_1__25_, nextQ_1__24_, 
        nextQ_1__23_, nextQ_1__22_, nextQ_1__21_, nextQ_1__20_, nextQ_1__19_, 
        nextQ_1__18_, nextQ_1__17_, nextQ_1__16_, nextQ_1__15_, nextQ_1__14_, 
        nextQ_1__13_, nextQ_1__12_, nextQ_1__11_, nextQ_1__10_, nextQ_1__9_, 
        nextQ_1__8_, nextQ_1__7_, nextQ_1__6_, nextQ_1__5_, nextQ_1__4_, 
        nextQ_1__3_, nextQ_1__2_, nextQ_1__1_, nextQ_1__0_}), .nextQ_1(q_1[1])
         );
  BoothStep_31 booth_instances_1__stepX ( .a({nextA_1__31_, nextA_1__30_, 
        nextA_1__29_, nextA_1__28_, nextA_1__27_, nextA_1__26_, nextA_1__25_, 
        nextA_1__24_, nextA_1__23_, nextA_1__22_, nextA_1__21_, nextA_1__20_, 
        nextA_1__19_, nextA_1__18_, nextA_1__17_, nextA_1__16_, nextA_1__15_, 
        nextA_1__14_, nextA_1__13_, nextA_1__12_, nextA_1__11_, nextA_1__10_, 
        nextA_1__9_, nextA_1__8_, nextA_1__7_, nextA_1__6_, nextA_1__5_, 
        nextA_1__4_, nextA_1__3_, nextA_1__2_, nextA_1__1_, nextA_1__0_}), .q(
        {nextQ_1__31_, nextQ_1__30_, nextQ_1__29_, nextQ_1__28_, nextQ_1__27_, 
        nextQ_1__26_, nextQ_1__25_, nextQ_1__24_, nextQ_1__23_, nextQ_1__22_, 
        nextQ_1__21_, nextQ_1__20_, nextQ_1__19_, nextQ_1__18_, nextQ_1__17_, 
        nextQ_1__16_, nextQ_1__15_, nextQ_1__14_, nextQ_1__13_, nextQ_1__12_, 
        nextQ_1__11_, nextQ_1__10_, nextQ_1__9_, nextQ_1__8_, nextQ_1__7_, 
        nextQ_1__6_, nextQ_1__5_, nextQ_1__4_, nextQ_1__3_, nextQ_1__2_, 
        nextQ_1__1_, nextQ_1__0_}), .m(a), .q_1(q_1[1]), .nextA({nextA_2__31_, 
        nextA_2__30_, nextA_2__29_, nextA_2__28_, nextA_2__27_, nextA_2__26_, 
        nextA_2__25_, nextA_2__24_, nextA_2__23_, nextA_2__22_, nextA_2__21_, 
        nextA_2__20_, nextA_2__19_, nextA_2__18_, nextA_2__17_, nextA_2__16_, 
        nextA_2__15_, nextA_2__14_, nextA_2__13_, nextA_2__12_, nextA_2__11_, 
        nextA_2__10_, nextA_2__9_, nextA_2__8_, nextA_2__7_, nextA_2__6_, 
        nextA_2__5_, nextA_2__4_, nextA_2__3_, nextA_2__2_, nextA_2__1_, 
        nextA_2__0_}), .nextQ({nextQ_2__31_, nextQ_2__30_, nextQ_2__29_, 
        nextQ_2__28_, nextQ_2__27_, nextQ_2__26_, nextQ_2__25_, nextQ_2__24_, 
        nextQ_2__23_, nextQ_2__22_, nextQ_2__21_, nextQ_2__20_, nextQ_2__19_, 
        nextQ_2__18_, nextQ_2__17_, nextQ_2__16_, nextQ_2__15_, nextQ_2__14_, 
        nextQ_2__13_, nextQ_2__12_, nextQ_2__11_, nextQ_2__10_, nextQ_2__9_, 
        nextQ_2__8_, nextQ_2__7_, nextQ_2__6_, nextQ_2__5_, nextQ_2__4_, 
        nextQ_2__3_, nextQ_2__2_, nextQ_2__1_, nextQ_2__0_}), .nextQ_1(q_1[2])
         );
  BoothStep_30 booth_instances_2__stepX ( .a({nextA_2__31_, nextA_2__30_, 
        nextA_2__29_, nextA_2__28_, nextA_2__27_, nextA_2__26_, nextA_2__25_, 
        nextA_2__24_, nextA_2__23_, nextA_2__22_, nextA_2__21_, nextA_2__20_, 
        nextA_2__19_, nextA_2__18_, nextA_2__17_, nextA_2__16_, nextA_2__15_, 
        nextA_2__14_, nextA_2__13_, nextA_2__12_, nextA_2__11_, nextA_2__10_, 
        nextA_2__9_, nextA_2__8_, nextA_2__7_, nextA_2__6_, nextA_2__5_, 
        nextA_2__4_, nextA_2__3_, nextA_2__2_, nextA_2__1_, nextA_2__0_}), .q(
        {nextQ_2__31_, nextQ_2__30_, nextQ_2__29_, nextQ_2__28_, nextQ_2__27_, 
        nextQ_2__26_, nextQ_2__25_, nextQ_2__24_, nextQ_2__23_, nextQ_2__22_, 
        nextQ_2__21_, nextQ_2__20_, nextQ_2__19_, nextQ_2__18_, nextQ_2__17_, 
        nextQ_2__16_, nextQ_2__15_, nextQ_2__14_, nextQ_2__13_, nextQ_2__12_, 
        nextQ_2__11_, nextQ_2__10_, nextQ_2__9_, nextQ_2__8_, nextQ_2__7_, 
        nextQ_2__6_, nextQ_2__5_, nextQ_2__4_, nextQ_2__3_, nextQ_2__2_, 
        nextQ_2__1_, nextQ_2__0_}), .m(a), .q_1(q_1[2]), .nextA({nextA_3__31_, 
        nextA_3__30_, nextA_3__29_, nextA_3__28_, nextA_3__27_, nextA_3__26_, 
        nextA_3__25_, nextA_3__24_, nextA_3__23_, nextA_3__22_, nextA_3__21_, 
        nextA_3__20_, nextA_3__19_, nextA_3__18_, nextA_3__17_, nextA_3__16_, 
        nextA_3__15_, nextA_3__14_, nextA_3__13_, nextA_3__12_, nextA_3__11_, 
        nextA_3__10_, nextA_3__9_, nextA_3__8_, nextA_3__7_, nextA_3__6_, 
        nextA_3__5_, nextA_3__4_, nextA_3__3_, nextA_3__2_, nextA_3__1_, 
        nextA_3__0_}), .nextQ({nextQ_3__31_, nextQ_3__30_, nextQ_3__29_, 
        nextQ_3__28_, nextQ_3__27_, nextQ_3__26_, nextQ_3__25_, nextQ_3__24_, 
        nextQ_3__23_, nextQ_3__22_, nextQ_3__21_, nextQ_3__20_, nextQ_3__19_, 
        nextQ_3__18_, nextQ_3__17_, nextQ_3__16_, nextQ_3__15_, nextQ_3__14_, 
        nextQ_3__13_, nextQ_3__12_, nextQ_3__11_, nextQ_3__10_, nextQ_3__9_, 
        nextQ_3__8_, nextQ_3__7_, nextQ_3__6_, nextQ_3__5_, nextQ_3__4_, 
        nextQ_3__3_, nextQ_3__2_, nextQ_3__1_, nextQ_3__0_}), .nextQ_1(q_1[3])
         );
  BoothStep_29 booth_instances_3__stepX ( .a({nextA_3__31_, nextA_3__30_, 
        nextA_3__29_, nextA_3__28_, nextA_3__27_, nextA_3__26_, nextA_3__25_, 
        nextA_3__24_, nextA_3__23_, nextA_3__22_, nextA_3__21_, nextA_3__20_, 
        nextA_3__19_, nextA_3__18_, nextA_3__17_, nextA_3__16_, nextA_3__15_, 
        nextA_3__14_, nextA_3__13_, nextA_3__12_, nextA_3__11_, nextA_3__10_, 
        nextA_3__9_, nextA_3__8_, nextA_3__7_, nextA_3__6_, nextA_3__5_, 
        nextA_3__4_, nextA_3__3_, nextA_3__2_, nextA_3__1_, nextA_3__0_}), .q(
        {nextQ_3__31_, nextQ_3__30_, nextQ_3__29_, nextQ_3__28_, nextQ_3__27_, 
        nextQ_3__26_, nextQ_3__25_, nextQ_3__24_, nextQ_3__23_, nextQ_3__22_, 
        nextQ_3__21_, nextQ_3__20_, nextQ_3__19_, nextQ_3__18_, nextQ_3__17_, 
        nextQ_3__16_, nextQ_3__15_, nextQ_3__14_, nextQ_3__13_, nextQ_3__12_, 
        nextQ_3__11_, nextQ_3__10_, nextQ_3__9_, nextQ_3__8_, nextQ_3__7_, 
        nextQ_3__6_, nextQ_3__5_, nextQ_3__4_, nextQ_3__3_, nextQ_3__2_, 
        nextQ_3__1_, nextQ_3__0_}), .m(a), .q_1(q_1[3]), .nextA({nextA_4__31_, 
        nextA_4__30_, nextA_4__29_, nextA_4__28_, nextA_4__27_, nextA_4__26_, 
        nextA_4__25_, nextA_4__24_, nextA_4__23_, nextA_4__22_, nextA_4__21_, 
        nextA_4__20_, nextA_4__19_, nextA_4__18_, nextA_4__17_, nextA_4__16_, 
        nextA_4__15_, nextA_4__14_, nextA_4__13_, nextA_4__12_, nextA_4__11_, 
        nextA_4__10_, nextA_4__9_, nextA_4__8_, nextA_4__7_, nextA_4__6_, 
        nextA_4__5_, nextA_4__4_, nextA_4__3_, nextA_4__2_, nextA_4__1_, 
        nextA_4__0_}), .nextQ({nextQ_4__31_, nextQ_4__30_, nextQ_4__29_, 
        nextQ_4__28_, nextQ_4__27_, nextQ_4__26_, nextQ_4__25_, nextQ_4__24_, 
        nextQ_4__23_, nextQ_4__22_, nextQ_4__21_, nextQ_4__20_, nextQ_4__19_, 
        nextQ_4__18_, nextQ_4__17_, nextQ_4__16_, nextQ_4__15_, nextQ_4__14_, 
        nextQ_4__13_, nextQ_4__12_, nextQ_4__11_, nextQ_4__10_, nextQ_4__9_, 
        nextQ_4__8_, nextQ_4__7_, nextQ_4__6_, nextQ_4__5_, nextQ_4__4_, 
        nextQ_4__3_, nextQ_4__2_, nextQ_4__1_, nextQ_4__0_}), .nextQ_1(q_1[4])
         );
  BoothStep_28 booth_instances_4__stepX ( .a({nextA_4__31_, nextA_4__30_, 
        nextA_4__29_, nextA_4__28_, nextA_4__27_, nextA_4__26_, nextA_4__25_, 
        nextA_4__24_, nextA_4__23_, nextA_4__22_, nextA_4__21_, nextA_4__20_, 
        nextA_4__19_, nextA_4__18_, nextA_4__17_, nextA_4__16_, nextA_4__15_, 
        nextA_4__14_, nextA_4__13_, nextA_4__12_, nextA_4__11_, nextA_4__10_, 
        nextA_4__9_, nextA_4__8_, nextA_4__7_, nextA_4__6_, nextA_4__5_, 
        nextA_4__4_, nextA_4__3_, nextA_4__2_, nextA_4__1_, nextA_4__0_}), .q(
        {nextQ_4__31_, nextQ_4__30_, nextQ_4__29_, nextQ_4__28_, nextQ_4__27_, 
        nextQ_4__26_, nextQ_4__25_, nextQ_4__24_, nextQ_4__23_, nextQ_4__22_, 
        nextQ_4__21_, nextQ_4__20_, nextQ_4__19_, nextQ_4__18_, nextQ_4__17_, 
        nextQ_4__16_, nextQ_4__15_, nextQ_4__14_, nextQ_4__13_, nextQ_4__12_, 
        nextQ_4__11_, nextQ_4__10_, nextQ_4__9_, nextQ_4__8_, nextQ_4__7_, 
        nextQ_4__6_, nextQ_4__5_, nextQ_4__4_, nextQ_4__3_, nextQ_4__2_, 
        nextQ_4__1_, nextQ_4__0_}), .m(a), .q_1(q_1[4]), .nextA({nextA_5__31_, 
        nextA_5__30_, nextA_5__29_, nextA_5__28_, nextA_5__27_, nextA_5__26_, 
        nextA_5__25_, nextA_5__24_, nextA_5__23_, nextA_5__22_, nextA_5__21_, 
        nextA_5__20_, nextA_5__19_, nextA_5__18_, nextA_5__17_, nextA_5__16_, 
        nextA_5__15_, nextA_5__14_, nextA_5__13_, nextA_5__12_, nextA_5__11_, 
        nextA_5__10_, nextA_5__9_, nextA_5__8_, nextA_5__7_, nextA_5__6_, 
        nextA_5__5_, nextA_5__4_, nextA_5__3_, nextA_5__2_, nextA_5__1_, 
        nextA_5__0_}), .nextQ({nextQ_5__31_, nextQ_5__30_, nextQ_5__29_, 
        nextQ_5__28_, nextQ_5__27_, nextQ_5__26_, nextQ_5__25_, nextQ_5__24_, 
        nextQ_5__23_, nextQ_5__22_, nextQ_5__21_, nextQ_5__20_, nextQ_5__19_, 
        nextQ_5__18_, nextQ_5__17_, nextQ_5__16_, nextQ_5__15_, nextQ_5__14_, 
        nextQ_5__13_, nextQ_5__12_, nextQ_5__11_, nextQ_5__10_, nextQ_5__9_, 
        nextQ_5__8_, nextQ_5__7_, nextQ_5__6_, nextQ_5__5_, nextQ_5__4_, 
        nextQ_5__3_, nextQ_5__2_, nextQ_5__1_, nextQ_5__0_}), .nextQ_1(q_1[5])
         );
  BoothStep_27 booth_instances_5__stepX ( .a({nextA_5__31_, nextA_5__30_, 
        nextA_5__29_, nextA_5__28_, nextA_5__27_, nextA_5__26_, nextA_5__25_, 
        nextA_5__24_, nextA_5__23_, nextA_5__22_, nextA_5__21_, nextA_5__20_, 
        nextA_5__19_, nextA_5__18_, nextA_5__17_, nextA_5__16_, nextA_5__15_, 
        nextA_5__14_, nextA_5__13_, nextA_5__12_, nextA_5__11_, nextA_5__10_, 
        nextA_5__9_, nextA_5__8_, nextA_5__7_, nextA_5__6_, nextA_5__5_, 
        nextA_5__4_, nextA_5__3_, nextA_5__2_, nextA_5__1_, nextA_5__0_}), .q(
        {nextQ_5__31_, nextQ_5__30_, nextQ_5__29_, nextQ_5__28_, nextQ_5__27_, 
        nextQ_5__26_, nextQ_5__25_, nextQ_5__24_, nextQ_5__23_, nextQ_5__22_, 
        nextQ_5__21_, nextQ_5__20_, nextQ_5__19_, nextQ_5__18_, nextQ_5__17_, 
        nextQ_5__16_, nextQ_5__15_, nextQ_5__14_, nextQ_5__13_, nextQ_5__12_, 
        nextQ_5__11_, nextQ_5__10_, nextQ_5__9_, nextQ_5__8_, nextQ_5__7_, 
        nextQ_5__6_, nextQ_5__5_, nextQ_5__4_, nextQ_5__3_, nextQ_5__2_, 
        nextQ_5__1_, nextQ_5__0_}), .m(a), .q_1(q_1[5]), .nextA({nextA_6__31_, 
        nextA_6__30_, nextA_6__29_, nextA_6__28_, nextA_6__27_, nextA_6__26_, 
        nextA_6__25_, nextA_6__24_, nextA_6__23_, nextA_6__22_, nextA_6__21_, 
        nextA_6__20_, nextA_6__19_, nextA_6__18_, nextA_6__17_, nextA_6__16_, 
        nextA_6__15_, nextA_6__14_, nextA_6__13_, nextA_6__12_, nextA_6__11_, 
        nextA_6__10_, nextA_6__9_, nextA_6__8_, nextA_6__7_, nextA_6__6_, 
        nextA_6__5_, nextA_6__4_, nextA_6__3_, nextA_6__2_, nextA_6__1_, 
        nextA_6__0_}), .nextQ({nextQ_6__31_, nextQ_6__30_, nextQ_6__29_, 
        nextQ_6__28_, nextQ_6__27_, nextQ_6__26_, nextQ_6__25_, nextQ_6__24_, 
        nextQ_6__23_, nextQ_6__22_, nextQ_6__21_, nextQ_6__20_, nextQ_6__19_, 
        nextQ_6__18_, nextQ_6__17_, nextQ_6__16_, nextQ_6__15_, nextQ_6__14_, 
        nextQ_6__13_, nextQ_6__12_, nextQ_6__11_, nextQ_6__10_, nextQ_6__9_, 
        nextQ_6__8_, nextQ_6__7_, nextQ_6__6_, nextQ_6__5_, nextQ_6__4_, 
        nextQ_6__3_, nextQ_6__2_, nextQ_6__1_, nextQ_6__0_}), .nextQ_1(q_1[6])
         );
  BoothStep_26 booth_instances_6__stepX ( .a({nextA_6__31_, nextA_6__30_, 
        nextA_6__29_, nextA_6__28_, nextA_6__27_, nextA_6__26_, nextA_6__25_, 
        nextA_6__24_, nextA_6__23_, nextA_6__22_, nextA_6__21_, nextA_6__20_, 
        nextA_6__19_, nextA_6__18_, nextA_6__17_, nextA_6__16_, nextA_6__15_, 
        nextA_6__14_, nextA_6__13_, nextA_6__12_, nextA_6__11_, nextA_6__10_, 
        nextA_6__9_, nextA_6__8_, nextA_6__7_, nextA_6__6_, nextA_6__5_, 
        nextA_6__4_, nextA_6__3_, nextA_6__2_, nextA_6__1_, nextA_6__0_}), .q(
        {nextQ_6__31_, nextQ_6__30_, nextQ_6__29_, nextQ_6__28_, nextQ_6__27_, 
        nextQ_6__26_, nextQ_6__25_, nextQ_6__24_, nextQ_6__23_, nextQ_6__22_, 
        nextQ_6__21_, nextQ_6__20_, nextQ_6__19_, nextQ_6__18_, nextQ_6__17_, 
        nextQ_6__16_, nextQ_6__15_, nextQ_6__14_, nextQ_6__13_, nextQ_6__12_, 
        nextQ_6__11_, nextQ_6__10_, nextQ_6__9_, nextQ_6__8_, nextQ_6__7_, 
        nextQ_6__6_, nextQ_6__5_, nextQ_6__4_, nextQ_6__3_, nextQ_6__2_, 
        nextQ_6__1_, nextQ_6__0_}), .m(a), .q_1(q_1[6]), .nextA({nextA_7__31_, 
        nextA_7__30_, nextA_7__29_, nextA_7__28_, nextA_7__27_, nextA_7__26_, 
        nextA_7__25_, nextA_7__24_, nextA_7__23_, nextA_7__22_, nextA_7__21_, 
        nextA_7__20_, nextA_7__19_, nextA_7__18_, nextA_7__17_, nextA_7__16_, 
        nextA_7__15_, nextA_7__14_, nextA_7__13_, nextA_7__12_, nextA_7__11_, 
        nextA_7__10_, nextA_7__9_, nextA_7__8_, nextA_7__7_, nextA_7__6_, 
        nextA_7__5_, nextA_7__4_, nextA_7__3_, nextA_7__2_, nextA_7__1_, 
        nextA_7__0_}), .nextQ({nextQ_7__31_, nextQ_7__30_, nextQ_7__29_, 
        nextQ_7__28_, nextQ_7__27_, nextQ_7__26_, nextQ_7__25_, nextQ_7__24_, 
        nextQ_7__23_, nextQ_7__22_, nextQ_7__21_, nextQ_7__20_, nextQ_7__19_, 
        nextQ_7__18_, nextQ_7__17_, nextQ_7__16_, nextQ_7__15_, nextQ_7__14_, 
        nextQ_7__13_, nextQ_7__12_, nextQ_7__11_, nextQ_7__10_, nextQ_7__9_, 
        nextQ_7__8_, nextQ_7__7_, nextQ_7__6_, nextQ_7__5_, nextQ_7__4_, 
        nextQ_7__3_, nextQ_7__2_, nextQ_7__1_, nextQ_7__0_}), .nextQ_1(q_1[7])
         );
  BoothStep_25 booth_instances_7__stepX ( .a({nextA_7__31_, nextA_7__30_, 
        nextA_7__29_, nextA_7__28_, nextA_7__27_, nextA_7__26_, nextA_7__25_, 
        nextA_7__24_, nextA_7__23_, nextA_7__22_, nextA_7__21_, nextA_7__20_, 
        nextA_7__19_, nextA_7__18_, nextA_7__17_, nextA_7__16_, nextA_7__15_, 
        nextA_7__14_, nextA_7__13_, nextA_7__12_, nextA_7__11_, nextA_7__10_, 
        nextA_7__9_, nextA_7__8_, nextA_7__7_, nextA_7__6_, nextA_7__5_, 
        nextA_7__4_, nextA_7__3_, nextA_7__2_, nextA_7__1_, nextA_7__0_}), .q(
        {nextQ_7__31_, nextQ_7__30_, nextQ_7__29_, nextQ_7__28_, nextQ_7__27_, 
        nextQ_7__26_, nextQ_7__25_, nextQ_7__24_, nextQ_7__23_, nextQ_7__22_, 
        nextQ_7__21_, nextQ_7__20_, nextQ_7__19_, nextQ_7__18_, nextQ_7__17_, 
        nextQ_7__16_, nextQ_7__15_, nextQ_7__14_, nextQ_7__13_, nextQ_7__12_, 
        nextQ_7__11_, nextQ_7__10_, nextQ_7__9_, nextQ_7__8_, nextQ_7__7_, 
        nextQ_7__6_, nextQ_7__5_, nextQ_7__4_, nextQ_7__3_, nextQ_7__2_, 
        nextQ_7__1_, nextQ_7__0_}), .m(a), .q_1(q_1[7]), .nextA({nextA_8__31_, 
        nextA_8__30_, nextA_8__29_, nextA_8__28_, nextA_8__27_, nextA_8__26_, 
        nextA_8__25_, nextA_8__24_, nextA_8__23_, nextA_8__22_, nextA_8__21_, 
        nextA_8__20_, nextA_8__19_, nextA_8__18_, nextA_8__17_, nextA_8__16_, 
        nextA_8__15_, nextA_8__14_, nextA_8__13_, nextA_8__12_, nextA_8__11_, 
        nextA_8__10_, nextA_8__9_, nextA_8__8_, nextA_8__7_, nextA_8__6_, 
        nextA_8__5_, nextA_8__4_, nextA_8__3_, nextA_8__2_, nextA_8__1_, 
        nextA_8__0_}), .nextQ({nextQ_8__31_, nextQ_8__30_, nextQ_8__29_, 
        nextQ_8__28_, nextQ_8__27_, nextQ_8__26_, nextQ_8__25_, nextQ_8__24_, 
        nextQ_8__23_, nextQ_8__22_, nextQ_8__21_, nextQ_8__20_, nextQ_8__19_, 
        nextQ_8__18_, nextQ_8__17_, nextQ_8__16_, nextQ_8__15_, nextQ_8__14_, 
        nextQ_8__13_, nextQ_8__12_, nextQ_8__11_, nextQ_8__10_, nextQ_8__9_, 
        nextQ_8__8_, nextQ_8__7_, nextQ_8__6_, nextQ_8__5_, nextQ_8__4_, 
        nextQ_8__3_, nextQ_8__2_, nextQ_8__1_, nextQ_8__0_}), .nextQ_1(q_1[8])
         );
  BoothStep_24 booth_instances_8__stepX ( .a({nextA_8__31_, nextA_8__30_, 
        nextA_8__29_, nextA_8__28_, nextA_8__27_, nextA_8__26_, nextA_8__25_, 
        nextA_8__24_, nextA_8__23_, nextA_8__22_, nextA_8__21_, nextA_8__20_, 
        nextA_8__19_, nextA_8__18_, nextA_8__17_, nextA_8__16_, nextA_8__15_, 
        nextA_8__14_, nextA_8__13_, nextA_8__12_, nextA_8__11_, nextA_8__10_, 
        nextA_8__9_, nextA_8__8_, nextA_8__7_, nextA_8__6_, nextA_8__5_, 
        nextA_8__4_, nextA_8__3_, nextA_8__2_, nextA_8__1_, nextA_8__0_}), .q(
        {nextQ_8__31_, nextQ_8__30_, nextQ_8__29_, nextQ_8__28_, nextQ_8__27_, 
        nextQ_8__26_, nextQ_8__25_, nextQ_8__24_, nextQ_8__23_, nextQ_8__22_, 
        nextQ_8__21_, nextQ_8__20_, nextQ_8__19_, nextQ_8__18_, nextQ_8__17_, 
        nextQ_8__16_, nextQ_8__15_, nextQ_8__14_, nextQ_8__13_, nextQ_8__12_, 
        nextQ_8__11_, nextQ_8__10_, nextQ_8__9_, nextQ_8__8_, nextQ_8__7_, 
        nextQ_8__6_, nextQ_8__5_, nextQ_8__4_, nextQ_8__3_, nextQ_8__2_, 
        nextQ_8__1_, nextQ_8__0_}), .m(a), .q_1(q_1[8]), .nextA({nextA_9__31_, 
        nextA_9__30_, nextA_9__29_, nextA_9__28_, nextA_9__27_, nextA_9__26_, 
        nextA_9__25_, nextA_9__24_, nextA_9__23_, nextA_9__22_, nextA_9__21_, 
        nextA_9__20_, nextA_9__19_, nextA_9__18_, nextA_9__17_, nextA_9__16_, 
        nextA_9__15_, nextA_9__14_, nextA_9__13_, nextA_9__12_, nextA_9__11_, 
        nextA_9__10_, nextA_9__9_, nextA_9__8_, nextA_9__7_, nextA_9__6_, 
        nextA_9__5_, nextA_9__4_, nextA_9__3_, nextA_9__2_, nextA_9__1_, 
        nextA_9__0_}), .nextQ({nextQ_9__31_, nextQ_9__30_, nextQ_9__29_, 
        nextQ_9__28_, nextQ_9__27_, nextQ_9__26_, nextQ_9__25_, nextQ_9__24_, 
        nextQ_9__23_, nextQ_9__22_, nextQ_9__21_, nextQ_9__20_, nextQ_9__19_, 
        nextQ_9__18_, nextQ_9__17_, nextQ_9__16_, nextQ_9__15_, nextQ_9__14_, 
        nextQ_9__13_, nextQ_9__12_, nextQ_9__11_, nextQ_9__10_, nextQ_9__9_, 
        nextQ_9__8_, nextQ_9__7_, nextQ_9__6_, nextQ_9__5_, nextQ_9__4_, 
        nextQ_9__3_, nextQ_9__2_, nextQ_9__1_, nextQ_9__0_}), .nextQ_1(q_1[9])
         );
  BoothStep_23 booth_instances_9__stepX ( .a({nextA_9__31_, nextA_9__30_, 
        nextA_9__29_, nextA_9__28_, nextA_9__27_, nextA_9__26_, nextA_9__25_, 
        nextA_9__24_, nextA_9__23_, nextA_9__22_, nextA_9__21_, nextA_9__20_, 
        nextA_9__19_, nextA_9__18_, nextA_9__17_, nextA_9__16_, nextA_9__15_, 
        nextA_9__14_, nextA_9__13_, nextA_9__12_, nextA_9__11_, nextA_9__10_, 
        nextA_9__9_, nextA_9__8_, nextA_9__7_, nextA_9__6_, nextA_9__5_, 
        nextA_9__4_, nextA_9__3_, nextA_9__2_, nextA_9__1_, nextA_9__0_}), .q(
        {nextQ_9__31_, nextQ_9__30_, nextQ_9__29_, nextQ_9__28_, nextQ_9__27_, 
        nextQ_9__26_, nextQ_9__25_, nextQ_9__24_, nextQ_9__23_, nextQ_9__22_, 
        nextQ_9__21_, nextQ_9__20_, nextQ_9__19_, nextQ_9__18_, nextQ_9__17_, 
        nextQ_9__16_, nextQ_9__15_, nextQ_9__14_, nextQ_9__13_, nextQ_9__12_, 
        nextQ_9__11_, nextQ_9__10_, nextQ_9__9_, nextQ_9__8_, nextQ_9__7_, 
        nextQ_9__6_, nextQ_9__5_, nextQ_9__4_, nextQ_9__3_, nextQ_9__2_, 
        nextQ_9__1_, nextQ_9__0_}), .m(a), .q_1(q_1[9]), .nextA({nextA_10__31_, 
        nextA_10__30_, nextA_10__29_, nextA_10__28_, nextA_10__27_, 
        nextA_10__26_, nextA_10__25_, nextA_10__24_, nextA_10__23_, 
        nextA_10__22_, nextA_10__21_, nextA_10__20_, nextA_10__19_, 
        nextA_10__18_, nextA_10__17_, nextA_10__16_, nextA_10__15_, 
        nextA_10__14_, nextA_10__13_, nextA_10__12_, nextA_10__11_, 
        nextA_10__10_, nextA_10__9_, nextA_10__8_, nextA_10__7_, nextA_10__6_, 
        nextA_10__5_, nextA_10__4_, nextA_10__3_, nextA_10__2_, nextA_10__1_, 
        nextA_10__0_}), .nextQ({nextQ_10__31_, nextQ_10__30_, nextQ_10__29_, 
        nextQ_10__28_, nextQ_10__27_, nextQ_10__26_, nextQ_10__25_, 
        nextQ_10__24_, nextQ_10__23_, nextQ_10__22_, nextQ_10__21_, 
        nextQ_10__20_, nextQ_10__19_, nextQ_10__18_, nextQ_10__17_, 
        nextQ_10__16_, nextQ_10__15_, nextQ_10__14_, nextQ_10__13_, 
        nextQ_10__12_, nextQ_10__11_, nextQ_10__10_, nextQ_10__9_, 
        nextQ_10__8_, nextQ_10__7_, nextQ_10__6_, nextQ_10__5_, nextQ_10__4_, 
        nextQ_10__3_, nextQ_10__2_, nextQ_10__1_, nextQ_10__0_}), .nextQ_1(
        q_1[10]) );
  BoothStep_22 booth_instances_10__stepX ( .a({nextA_10__31_, nextA_10__30_, 
        nextA_10__29_, nextA_10__28_, nextA_10__27_, nextA_10__26_, 
        nextA_10__25_, nextA_10__24_, nextA_10__23_, nextA_10__22_, 
        nextA_10__21_, nextA_10__20_, nextA_10__19_, nextA_10__18_, 
        nextA_10__17_, nextA_10__16_, nextA_10__15_, nextA_10__14_, 
        nextA_10__13_, nextA_10__12_, nextA_10__11_, nextA_10__10_, 
        nextA_10__9_, nextA_10__8_, nextA_10__7_, nextA_10__6_, nextA_10__5_, 
        nextA_10__4_, nextA_10__3_, nextA_10__2_, nextA_10__1_, nextA_10__0_}), 
        .q({nextQ_10__31_, nextQ_10__30_, nextQ_10__29_, nextQ_10__28_, 
        nextQ_10__27_, nextQ_10__26_, nextQ_10__25_, nextQ_10__24_, 
        nextQ_10__23_, nextQ_10__22_, nextQ_10__21_, nextQ_10__20_, 
        nextQ_10__19_, nextQ_10__18_, nextQ_10__17_, nextQ_10__16_, 
        nextQ_10__15_, nextQ_10__14_, nextQ_10__13_, nextQ_10__12_, 
        nextQ_10__11_, nextQ_10__10_, nextQ_10__9_, nextQ_10__8_, nextQ_10__7_, 
        nextQ_10__6_, nextQ_10__5_, nextQ_10__4_, nextQ_10__3_, nextQ_10__2_, 
        nextQ_10__1_, nextQ_10__0_}), .m(a), .q_1(q_1[10]), .nextA({
        nextA_11__31_, nextA_11__30_, nextA_11__29_, nextA_11__28_, 
        nextA_11__27_, nextA_11__26_, nextA_11__25_, nextA_11__24_, 
        nextA_11__23_, nextA_11__22_, nextA_11__21_, nextA_11__20_, 
        nextA_11__19_, nextA_11__18_, nextA_11__17_, nextA_11__16_, 
        nextA_11__15_, nextA_11__14_, nextA_11__13_, nextA_11__12_, 
        nextA_11__11_, nextA_11__10_, nextA_11__9_, nextA_11__8_, nextA_11__7_, 
        nextA_11__6_, nextA_11__5_, nextA_11__4_, nextA_11__3_, nextA_11__2_, 
        nextA_11__1_, nextA_11__0_}), .nextQ({nextQ_11__31_, nextQ_11__30_, 
        nextQ_11__29_, nextQ_11__28_, nextQ_11__27_, nextQ_11__26_, 
        nextQ_11__25_, nextQ_11__24_, nextQ_11__23_, nextQ_11__22_, 
        nextQ_11__21_, nextQ_11__20_, nextQ_11__19_, nextQ_11__18_, 
        nextQ_11__17_, nextQ_11__16_, nextQ_11__15_, nextQ_11__14_, 
        nextQ_11__13_, nextQ_11__12_, nextQ_11__11_, nextQ_11__10_, 
        nextQ_11__9_, nextQ_11__8_, nextQ_11__7_, nextQ_11__6_, nextQ_11__5_, 
        nextQ_11__4_, nextQ_11__3_, nextQ_11__2_, nextQ_11__1_, nextQ_11__0_}), 
        .nextQ_1(q_1[11]) );
  BoothStep_21 booth_instances_11__stepX ( .a({nextA_11__31_, nextA_11__30_, 
        nextA_11__29_, nextA_11__28_, nextA_11__27_, nextA_11__26_, 
        nextA_11__25_, nextA_11__24_, nextA_11__23_, nextA_11__22_, 
        nextA_11__21_, nextA_11__20_, nextA_11__19_, nextA_11__18_, 
        nextA_11__17_, nextA_11__16_, nextA_11__15_, nextA_11__14_, 
        nextA_11__13_, nextA_11__12_, nextA_11__11_, nextA_11__10_, 
        nextA_11__9_, nextA_11__8_, nextA_11__7_, nextA_11__6_, nextA_11__5_, 
        nextA_11__4_, nextA_11__3_, nextA_11__2_, nextA_11__1_, nextA_11__0_}), 
        .q({nextQ_11__31_, nextQ_11__30_, nextQ_11__29_, nextQ_11__28_, 
        nextQ_11__27_, nextQ_11__26_, nextQ_11__25_, nextQ_11__24_, 
        nextQ_11__23_, nextQ_11__22_, nextQ_11__21_, nextQ_11__20_, 
        nextQ_11__19_, nextQ_11__18_, nextQ_11__17_, nextQ_11__16_, 
        nextQ_11__15_, nextQ_11__14_, nextQ_11__13_, nextQ_11__12_, 
        nextQ_11__11_, nextQ_11__10_, nextQ_11__9_, nextQ_11__8_, nextQ_11__7_, 
        nextQ_11__6_, nextQ_11__5_, nextQ_11__4_, nextQ_11__3_, nextQ_11__2_, 
        nextQ_11__1_, nextQ_11__0_}), .m(a), .q_1(q_1[11]), .nextA({
        nextA_12__31_, nextA_12__30_, nextA_12__29_, nextA_12__28_, 
        nextA_12__27_, nextA_12__26_, nextA_12__25_, nextA_12__24_, 
        nextA_12__23_, nextA_12__22_, nextA_12__21_, nextA_12__20_, 
        nextA_12__19_, nextA_12__18_, nextA_12__17_, nextA_12__16_, 
        nextA_12__15_, nextA_12__14_, nextA_12__13_, nextA_12__12_, 
        nextA_12__11_, nextA_12__10_, nextA_12__9_, nextA_12__8_, nextA_12__7_, 
        nextA_12__6_, nextA_12__5_, nextA_12__4_, nextA_12__3_, nextA_12__2_, 
        nextA_12__1_, nextA_12__0_}), .nextQ({nextQ_12__31_, nextQ_12__30_, 
        nextQ_12__29_, nextQ_12__28_, nextQ_12__27_, nextQ_12__26_, 
        nextQ_12__25_, nextQ_12__24_, nextQ_12__23_, nextQ_12__22_, 
        nextQ_12__21_, nextQ_12__20_, nextQ_12__19_, nextQ_12__18_, 
        nextQ_12__17_, nextQ_12__16_, nextQ_12__15_, nextQ_12__14_, 
        nextQ_12__13_, nextQ_12__12_, nextQ_12__11_, nextQ_12__10_, 
        nextQ_12__9_, nextQ_12__8_, nextQ_12__7_, nextQ_12__6_, nextQ_12__5_, 
        nextQ_12__4_, nextQ_12__3_, nextQ_12__2_, nextQ_12__1_, nextQ_12__0_}), 
        .nextQ_1(q_1[12]) );
  BoothStep_20 booth_instances_12__stepX ( .a({nextA_12__31_, nextA_12__30_, 
        nextA_12__29_, nextA_12__28_, nextA_12__27_, nextA_12__26_, 
        nextA_12__25_, nextA_12__24_, nextA_12__23_, nextA_12__22_, 
        nextA_12__21_, nextA_12__20_, nextA_12__19_, nextA_12__18_, 
        nextA_12__17_, nextA_12__16_, nextA_12__15_, nextA_12__14_, 
        nextA_12__13_, nextA_12__12_, nextA_12__11_, nextA_12__10_, 
        nextA_12__9_, nextA_12__8_, nextA_12__7_, nextA_12__6_, nextA_12__5_, 
        nextA_12__4_, nextA_12__3_, nextA_12__2_, nextA_12__1_, nextA_12__0_}), 
        .q({nextQ_12__31_, nextQ_12__30_, nextQ_12__29_, nextQ_12__28_, 
        nextQ_12__27_, nextQ_12__26_, nextQ_12__25_, nextQ_12__24_, 
        nextQ_12__23_, nextQ_12__22_, nextQ_12__21_, nextQ_12__20_, 
        nextQ_12__19_, nextQ_12__18_, nextQ_12__17_, nextQ_12__16_, 
        nextQ_12__15_, nextQ_12__14_, nextQ_12__13_, nextQ_12__12_, 
        nextQ_12__11_, nextQ_12__10_, nextQ_12__9_, nextQ_12__8_, nextQ_12__7_, 
        nextQ_12__6_, nextQ_12__5_, nextQ_12__4_, nextQ_12__3_, nextQ_12__2_, 
        nextQ_12__1_, nextQ_12__0_}), .m(a), .q_1(q_1[12]), .nextA({
        nextA_13__31_, nextA_13__30_, nextA_13__29_, nextA_13__28_, 
        nextA_13__27_, nextA_13__26_, nextA_13__25_, nextA_13__24_, 
        nextA_13__23_, nextA_13__22_, nextA_13__21_, nextA_13__20_, 
        nextA_13__19_, nextA_13__18_, nextA_13__17_, nextA_13__16_, 
        nextA_13__15_, nextA_13__14_, nextA_13__13_, nextA_13__12_, 
        nextA_13__11_, nextA_13__10_, nextA_13__9_, nextA_13__8_, nextA_13__7_, 
        nextA_13__6_, nextA_13__5_, nextA_13__4_, nextA_13__3_, nextA_13__2_, 
        nextA_13__1_, nextA_13__0_}), .nextQ({nextQ_13__31_, nextQ_13__30_, 
        nextQ_13__29_, nextQ_13__28_, nextQ_13__27_, nextQ_13__26_, 
        nextQ_13__25_, nextQ_13__24_, nextQ_13__23_, nextQ_13__22_, 
        nextQ_13__21_, nextQ_13__20_, nextQ_13__19_, nextQ_13__18_, 
        nextQ_13__17_, nextQ_13__16_, nextQ_13__15_, nextQ_13__14_, 
        nextQ_13__13_, nextQ_13__12_, nextQ_13__11_, nextQ_13__10_, 
        nextQ_13__9_, nextQ_13__8_, nextQ_13__7_, nextQ_13__6_, nextQ_13__5_, 
        nextQ_13__4_, nextQ_13__3_, nextQ_13__2_, nextQ_13__1_, nextQ_13__0_}), 
        .nextQ_1(q_1[13]) );
  BoothStep_19 booth_instances_13__stepX ( .a({nextA_13__31_, nextA_13__30_, 
        nextA_13__29_, nextA_13__28_, nextA_13__27_, nextA_13__26_, 
        nextA_13__25_, nextA_13__24_, nextA_13__23_, nextA_13__22_, 
        nextA_13__21_, nextA_13__20_, nextA_13__19_, nextA_13__18_, 
        nextA_13__17_, nextA_13__16_, nextA_13__15_, nextA_13__14_, 
        nextA_13__13_, nextA_13__12_, nextA_13__11_, nextA_13__10_, 
        nextA_13__9_, nextA_13__8_, nextA_13__7_, nextA_13__6_, nextA_13__5_, 
        nextA_13__4_, nextA_13__3_, nextA_13__2_, nextA_13__1_, nextA_13__0_}), 
        .q({nextQ_13__31_, nextQ_13__30_, nextQ_13__29_, nextQ_13__28_, 
        nextQ_13__27_, nextQ_13__26_, nextQ_13__25_, nextQ_13__24_, 
        nextQ_13__23_, nextQ_13__22_, nextQ_13__21_, nextQ_13__20_, 
        nextQ_13__19_, nextQ_13__18_, nextQ_13__17_, nextQ_13__16_, 
        nextQ_13__15_, nextQ_13__14_, nextQ_13__13_, nextQ_13__12_, 
        nextQ_13__11_, nextQ_13__10_, nextQ_13__9_, nextQ_13__8_, nextQ_13__7_, 
        nextQ_13__6_, nextQ_13__5_, nextQ_13__4_, nextQ_13__3_, nextQ_13__2_, 
        nextQ_13__1_, nextQ_13__0_}), .m(a), .q_1(q_1[13]), .nextA({
        nextA_14__31_, nextA_14__30_, nextA_14__29_, nextA_14__28_, 
        nextA_14__27_, nextA_14__26_, nextA_14__25_, nextA_14__24_, 
        nextA_14__23_, nextA_14__22_, nextA_14__21_, nextA_14__20_, 
        nextA_14__19_, nextA_14__18_, nextA_14__17_, nextA_14__16_, 
        nextA_14__15_, nextA_14__14_, nextA_14__13_, nextA_14__12_, 
        nextA_14__11_, nextA_14__10_, nextA_14__9_, nextA_14__8_, nextA_14__7_, 
        nextA_14__6_, nextA_14__5_, nextA_14__4_, nextA_14__3_, nextA_14__2_, 
        nextA_14__1_, nextA_14__0_}), .nextQ({nextQ_14__31_, nextQ_14__30_, 
        nextQ_14__29_, nextQ_14__28_, nextQ_14__27_, nextQ_14__26_, 
        nextQ_14__25_, nextQ_14__24_, nextQ_14__23_, nextQ_14__22_, 
        nextQ_14__21_, nextQ_14__20_, nextQ_14__19_, nextQ_14__18_, 
        nextQ_14__17_, nextQ_14__16_, nextQ_14__15_, nextQ_14__14_, 
        nextQ_14__13_, nextQ_14__12_, nextQ_14__11_, nextQ_14__10_, 
        nextQ_14__9_, nextQ_14__8_, nextQ_14__7_, nextQ_14__6_, nextQ_14__5_, 
        nextQ_14__4_, nextQ_14__3_, nextQ_14__2_, nextQ_14__1_, nextQ_14__0_}), 
        .nextQ_1(q_1[14]) );
  BoothStep_18 booth_instances_14__stepX ( .a({nextA_14__31_, nextA_14__30_, 
        nextA_14__29_, nextA_14__28_, nextA_14__27_, nextA_14__26_, 
        nextA_14__25_, nextA_14__24_, nextA_14__23_, nextA_14__22_, 
        nextA_14__21_, nextA_14__20_, nextA_14__19_, nextA_14__18_, 
        nextA_14__17_, nextA_14__16_, nextA_14__15_, nextA_14__14_, 
        nextA_14__13_, nextA_14__12_, nextA_14__11_, nextA_14__10_, 
        nextA_14__9_, nextA_14__8_, nextA_14__7_, nextA_14__6_, nextA_14__5_, 
        nextA_14__4_, nextA_14__3_, nextA_14__2_, nextA_14__1_, nextA_14__0_}), 
        .q({nextQ_14__31_, nextQ_14__30_, nextQ_14__29_, nextQ_14__28_, 
        nextQ_14__27_, nextQ_14__26_, nextQ_14__25_, nextQ_14__24_, 
        nextQ_14__23_, nextQ_14__22_, nextQ_14__21_, nextQ_14__20_, 
        nextQ_14__19_, nextQ_14__18_, nextQ_14__17_, nextQ_14__16_, 
        nextQ_14__15_, nextQ_14__14_, nextQ_14__13_, nextQ_14__12_, 
        nextQ_14__11_, nextQ_14__10_, nextQ_14__9_, nextQ_14__8_, nextQ_14__7_, 
        nextQ_14__6_, nextQ_14__5_, nextQ_14__4_, nextQ_14__3_, nextQ_14__2_, 
        nextQ_14__1_, nextQ_14__0_}), .m(a), .q_1(q_1[14]), .nextA({
        nextA_15__31_, nextA_15__30_, nextA_15__29_, nextA_15__28_, 
        nextA_15__27_, nextA_15__26_, nextA_15__25_, nextA_15__24_, 
        nextA_15__23_, nextA_15__22_, nextA_15__21_, nextA_15__20_, 
        nextA_15__19_, nextA_15__18_, nextA_15__17_, nextA_15__16_, 
        nextA_15__15_, nextA_15__14_, nextA_15__13_, nextA_15__12_, 
        nextA_15__11_, nextA_15__10_, nextA_15__9_, nextA_15__8_, nextA_15__7_, 
        nextA_15__6_, nextA_15__5_, nextA_15__4_, nextA_15__3_, nextA_15__2_, 
        nextA_15__1_, nextA_15__0_}), .nextQ({nextQ_15__31_, nextQ_15__30_, 
        nextQ_15__29_, nextQ_15__28_, nextQ_15__27_, nextQ_15__26_, 
        nextQ_15__25_, nextQ_15__24_, nextQ_15__23_, nextQ_15__22_, 
        nextQ_15__21_, nextQ_15__20_, nextQ_15__19_, nextQ_15__18_, 
        nextQ_15__17_, nextQ_15__16_, nextQ_15__15_, nextQ_15__14_, 
        nextQ_15__13_, nextQ_15__12_, nextQ_15__11_, nextQ_15__10_, 
        nextQ_15__9_, nextQ_15__8_, nextQ_15__7_, nextQ_15__6_, nextQ_15__5_, 
        nextQ_15__4_, nextQ_15__3_, nextQ_15__2_, nextQ_15__1_, nextQ_15__0_}), 
        .nextQ_1(q_1[15]) );
  BoothStep_17 booth_instances_15__stepX ( .a({nextA_15__31_, nextA_15__30_, 
        nextA_15__29_, nextA_15__28_, nextA_15__27_, nextA_15__26_, 
        nextA_15__25_, nextA_15__24_, nextA_15__23_, nextA_15__22_, 
        nextA_15__21_, nextA_15__20_, nextA_15__19_, nextA_15__18_, 
        nextA_15__17_, nextA_15__16_, nextA_15__15_, nextA_15__14_, 
        nextA_15__13_, nextA_15__12_, nextA_15__11_, nextA_15__10_, 
        nextA_15__9_, nextA_15__8_, nextA_15__7_, nextA_15__6_, nextA_15__5_, 
        nextA_15__4_, nextA_15__3_, nextA_15__2_, nextA_15__1_, nextA_15__0_}), 
        .q({nextQ_15__31_, nextQ_15__30_, nextQ_15__29_, nextQ_15__28_, 
        nextQ_15__27_, nextQ_15__26_, nextQ_15__25_, nextQ_15__24_, 
        nextQ_15__23_, nextQ_15__22_, nextQ_15__21_, nextQ_15__20_, 
        nextQ_15__19_, nextQ_15__18_, nextQ_15__17_, nextQ_15__16_, 
        nextQ_15__15_, nextQ_15__14_, nextQ_15__13_, nextQ_15__12_, 
        nextQ_15__11_, nextQ_15__10_, nextQ_15__9_, nextQ_15__8_, nextQ_15__7_, 
        nextQ_15__6_, nextQ_15__5_, nextQ_15__4_, nextQ_15__3_, nextQ_15__2_, 
        nextQ_15__1_, nextQ_15__0_}), .m(a), .q_1(q_1[15]), .nextA({
        nextA_16__31_, nextA_16__30_, nextA_16__29_, nextA_16__28_, 
        nextA_16__27_, nextA_16__26_, nextA_16__25_, nextA_16__24_, 
        nextA_16__23_, nextA_16__22_, nextA_16__21_, nextA_16__20_, 
        nextA_16__19_, nextA_16__18_, nextA_16__17_, nextA_16__16_, 
        nextA_16__15_, nextA_16__14_, nextA_16__13_, nextA_16__12_, 
        nextA_16__11_, nextA_16__10_, nextA_16__9_, nextA_16__8_, nextA_16__7_, 
        nextA_16__6_, nextA_16__5_, nextA_16__4_, nextA_16__3_, nextA_16__2_, 
        nextA_16__1_, nextA_16__0_}), .nextQ({nextQ_16__31_, nextQ_16__30_, 
        nextQ_16__29_, nextQ_16__28_, nextQ_16__27_, nextQ_16__26_, 
        nextQ_16__25_, nextQ_16__24_, nextQ_16__23_, nextQ_16__22_, 
        nextQ_16__21_, nextQ_16__20_, nextQ_16__19_, nextQ_16__18_, 
        nextQ_16__17_, nextQ_16__16_, nextQ_16__15_, nextQ_16__14_, 
        nextQ_16__13_, nextQ_16__12_, nextQ_16__11_, nextQ_16__10_, 
        nextQ_16__9_, nextQ_16__8_, nextQ_16__7_, nextQ_16__6_, nextQ_16__5_, 
        nextQ_16__4_, nextQ_16__3_, nextQ_16__2_, nextQ_16__1_, nextQ_16__0_}), 
        .nextQ_1(q_1[16]) );
  BoothStep_16 booth_instances_16__stepX ( .a({nextA_16__31_, nextA_16__30_, 
        nextA_16__29_, nextA_16__28_, nextA_16__27_, nextA_16__26_, 
        nextA_16__25_, nextA_16__24_, nextA_16__23_, nextA_16__22_, 
        nextA_16__21_, nextA_16__20_, nextA_16__19_, nextA_16__18_, 
        nextA_16__17_, nextA_16__16_, nextA_16__15_, nextA_16__14_, 
        nextA_16__13_, nextA_16__12_, nextA_16__11_, nextA_16__10_, 
        nextA_16__9_, nextA_16__8_, nextA_16__7_, nextA_16__6_, nextA_16__5_, 
        nextA_16__4_, nextA_16__3_, nextA_16__2_, nextA_16__1_, nextA_16__0_}), 
        .q({nextQ_16__31_, nextQ_16__30_, nextQ_16__29_, nextQ_16__28_, 
        nextQ_16__27_, nextQ_16__26_, nextQ_16__25_, nextQ_16__24_, 
        nextQ_16__23_, nextQ_16__22_, nextQ_16__21_, nextQ_16__20_, 
        nextQ_16__19_, nextQ_16__18_, nextQ_16__17_, nextQ_16__16_, 
        nextQ_16__15_, nextQ_16__14_, nextQ_16__13_, nextQ_16__12_, 
        nextQ_16__11_, nextQ_16__10_, nextQ_16__9_, nextQ_16__8_, nextQ_16__7_, 
        nextQ_16__6_, nextQ_16__5_, nextQ_16__4_, nextQ_16__3_, nextQ_16__2_, 
        nextQ_16__1_, nextQ_16__0_}), .m(a), .q_1(q_1[16]), .nextA({
        nextA_17__31_, nextA_17__30_, nextA_17__29_, nextA_17__28_, 
        nextA_17__27_, nextA_17__26_, nextA_17__25_, nextA_17__24_, 
        nextA_17__23_, nextA_17__22_, nextA_17__21_, nextA_17__20_, 
        nextA_17__19_, nextA_17__18_, nextA_17__17_, nextA_17__16_, 
        nextA_17__15_, nextA_17__14_, nextA_17__13_, nextA_17__12_, 
        nextA_17__11_, nextA_17__10_, nextA_17__9_, nextA_17__8_, nextA_17__7_, 
        nextA_17__6_, nextA_17__5_, nextA_17__4_, nextA_17__3_, nextA_17__2_, 
        nextA_17__1_, nextA_17__0_}), .nextQ({nextQ_17__31_, nextQ_17__30_, 
        nextQ_17__29_, nextQ_17__28_, nextQ_17__27_, nextQ_17__26_, 
        nextQ_17__25_, nextQ_17__24_, nextQ_17__23_, nextQ_17__22_, 
        nextQ_17__21_, nextQ_17__20_, nextQ_17__19_, nextQ_17__18_, 
        nextQ_17__17_, nextQ_17__16_, nextQ_17__15_, nextQ_17__14_, 
        nextQ_17__13_, nextQ_17__12_, nextQ_17__11_, nextQ_17__10_, 
        nextQ_17__9_, nextQ_17__8_, nextQ_17__7_, nextQ_17__6_, nextQ_17__5_, 
        nextQ_17__4_, nextQ_17__3_, nextQ_17__2_, nextQ_17__1_, nextQ_17__0_}), 
        .nextQ_1(q_1[17]) );
  BoothStep_15 booth_instances_17__stepX ( .a({nextA_17__31_, nextA_17__30_, 
        nextA_17__29_, nextA_17__28_, nextA_17__27_, nextA_17__26_, 
        nextA_17__25_, nextA_17__24_, nextA_17__23_, nextA_17__22_, 
        nextA_17__21_, nextA_17__20_, nextA_17__19_, nextA_17__18_, 
        nextA_17__17_, nextA_17__16_, nextA_17__15_, nextA_17__14_, 
        nextA_17__13_, nextA_17__12_, nextA_17__11_, nextA_17__10_, 
        nextA_17__9_, nextA_17__8_, nextA_17__7_, nextA_17__6_, nextA_17__5_, 
        nextA_17__4_, nextA_17__3_, nextA_17__2_, nextA_17__1_, nextA_17__0_}), 
        .q({nextQ_17__31_, nextQ_17__30_, nextQ_17__29_, nextQ_17__28_, 
        nextQ_17__27_, nextQ_17__26_, nextQ_17__25_, nextQ_17__24_, 
        nextQ_17__23_, nextQ_17__22_, nextQ_17__21_, nextQ_17__20_, 
        nextQ_17__19_, nextQ_17__18_, nextQ_17__17_, nextQ_17__16_, 
        nextQ_17__15_, nextQ_17__14_, nextQ_17__13_, nextQ_17__12_, 
        nextQ_17__11_, nextQ_17__10_, nextQ_17__9_, nextQ_17__8_, nextQ_17__7_, 
        nextQ_17__6_, nextQ_17__5_, nextQ_17__4_, nextQ_17__3_, nextQ_17__2_, 
        nextQ_17__1_, nextQ_17__0_}), .m(a), .q_1(q_1[17]), .nextA({
        nextA_18__31_, nextA_18__30_, nextA_18__29_, nextA_18__28_, 
        nextA_18__27_, nextA_18__26_, nextA_18__25_, nextA_18__24_, 
        nextA_18__23_, nextA_18__22_, nextA_18__21_, nextA_18__20_, 
        nextA_18__19_, nextA_18__18_, nextA_18__17_, nextA_18__16_, 
        nextA_18__15_, nextA_18__14_, nextA_18__13_, nextA_18__12_, 
        nextA_18__11_, nextA_18__10_, nextA_18__9_, nextA_18__8_, nextA_18__7_, 
        nextA_18__6_, nextA_18__5_, nextA_18__4_, nextA_18__3_, nextA_18__2_, 
        nextA_18__1_, nextA_18__0_}), .nextQ({nextQ_18__31_, nextQ_18__30_, 
        nextQ_18__29_, nextQ_18__28_, nextQ_18__27_, nextQ_18__26_, 
        nextQ_18__25_, nextQ_18__24_, nextQ_18__23_, nextQ_18__22_, 
        nextQ_18__21_, nextQ_18__20_, nextQ_18__19_, nextQ_18__18_, 
        nextQ_18__17_, nextQ_18__16_, nextQ_18__15_, nextQ_18__14_, 
        nextQ_18__13_, nextQ_18__12_, nextQ_18__11_, nextQ_18__10_, 
        nextQ_18__9_, nextQ_18__8_, nextQ_18__7_, nextQ_18__6_, nextQ_18__5_, 
        nextQ_18__4_, nextQ_18__3_, nextQ_18__2_, nextQ_18__1_, nextQ_18__0_}), 
        .nextQ_1(q_1[18]) );
  BoothStep_14 booth_instances_18__stepX ( .a({nextA_18__31_, nextA_18__30_, 
        nextA_18__29_, nextA_18__28_, nextA_18__27_, nextA_18__26_, 
        nextA_18__25_, nextA_18__24_, nextA_18__23_, nextA_18__22_, 
        nextA_18__21_, nextA_18__20_, nextA_18__19_, nextA_18__18_, 
        nextA_18__17_, nextA_18__16_, nextA_18__15_, nextA_18__14_, 
        nextA_18__13_, nextA_18__12_, nextA_18__11_, nextA_18__10_, 
        nextA_18__9_, nextA_18__8_, nextA_18__7_, nextA_18__6_, nextA_18__5_, 
        nextA_18__4_, nextA_18__3_, nextA_18__2_, nextA_18__1_, nextA_18__0_}), 
        .q({nextQ_18__31_, nextQ_18__30_, nextQ_18__29_, nextQ_18__28_, 
        nextQ_18__27_, nextQ_18__26_, nextQ_18__25_, nextQ_18__24_, 
        nextQ_18__23_, nextQ_18__22_, nextQ_18__21_, nextQ_18__20_, 
        nextQ_18__19_, nextQ_18__18_, nextQ_18__17_, nextQ_18__16_, 
        nextQ_18__15_, nextQ_18__14_, nextQ_18__13_, nextQ_18__12_, 
        nextQ_18__11_, nextQ_18__10_, nextQ_18__9_, nextQ_18__8_, nextQ_18__7_, 
        nextQ_18__6_, nextQ_18__5_, nextQ_18__4_, nextQ_18__3_, nextQ_18__2_, 
        nextQ_18__1_, nextQ_18__0_}), .m(a), .q_1(q_1[18]), .nextA({
        nextA_19__31_, nextA_19__30_, nextA_19__29_, nextA_19__28_, 
        nextA_19__27_, nextA_19__26_, nextA_19__25_, nextA_19__24_, 
        nextA_19__23_, nextA_19__22_, nextA_19__21_, nextA_19__20_, 
        nextA_19__19_, nextA_19__18_, nextA_19__17_, nextA_19__16_, 
        nextA_19__15_, nextA_19__14_, nextA_19__13_, nextA_19__12_, 
        nextA_19__11_, nextA_19__10_, nextA_19__9_, nextA_19__8_, nextA_19__7_, 
        nextA_19__6_, nextA_19__5_, nextA_19__4_, nextA_19__3_, nextA_19__2_, 
        nextA_19__1_, nextA_19__0_}), .nextQ({nextQ_19__31_, nextQ_19__30_, 
        nextQ_19__29_, nextQ_19__28_, nextQ_19__27_, nextQ_19__26_, 
        nextQ_19__25_, nextQ_19__24_, nextQ_19__23_, nextQ_19__22_, 
        nextQ_19__21_, nextQ_19__20_, nextQ_19__19_, nextQ_19__18_, 
        nextQ_19__17_, nextQ_19__16_, nextQ_19__15_, nextQ_19__14_, 
        nextQ_19__13_, nextQ_19__12_, nextQ_19__11_, nextQ_19__10_, 
        nextQ_19__9_, nextQ_19__8_, nextQ_19__7_, nextQ_19__6_, nextQ_19__5_, 
        nextQ_19__4_, nextQ_19__3_, nextQ_19__2_, nextQ_19__1_, nextQ_19__0_}), 
        .nextQ_1(q_1[19]) );
  BoothStep_13 booth_instances_19__stepX ( .a({nextA_19__31_, nextA_19__30_, 
        nextA_19__29_, nextA_19__28_, nextA_19__27_, nextA_19__26_, 
        nextA_19__25_, nextA_19__24_, nextA_19__23_, nextA_19__22_, 
        nextA_19__21_, nextA_19__20_, nextA_19__19_, nextA_19__18_, 
        nextA_19__17_, nextA_19__16_, nextA_19__15_, nextA_19__14_, 
        nextA_19__13_, nextA_19__12_, nextA_19__11_, nextA_19__10_, 
        nextA_19__9_, nextA_19__8_, nextA_19__7_, nextA_19__6_, nextA_19__5_, 
        nextA_19__4_, nextA_19__3_, nextA_19__2_, nextA_19__1_, nextA_19__0_}), 
        .q({nextQ_19__31_, nextQ_19__30_, nextQ_19__29_, nextQ_19__28_, 
        nextQ_19__27_, nextQ_19__26_, nextQ_19__25_, nextQ_19__24_, 
        nextQ_19__23_, nextQ_19__22_, nextQ_19__21_, nextQ_19__20_, 
        nextQ_19__19_, nextQ_19__18_, nextQ_19__17_, nextQ_19__16_, 
        nextQ_19__15_, nextQ_19__14_, nextQ_19__13_, nextQ_19__12_, 
        nextQ_19__11_, nextQ_19__10_, nextQ_19__9_, nextQ_19__8_, nextQ_19__7_, 
        nextQ_19__6_, nextQ_19__5_, nextQ_19__4_, nextQ_19__3_, nextQ_19__2_, 
        nextQ_19__1_, nextQ_19__0_}), .m(a), .q_1(q_1[19]), .nextA({
        nextA_20__31_, nextA_20__30_, nextA_20__29_, nextA_20__28_, 
        nextA_20__27_, nextA_20__26_, nextA_20__25_, nextA_20__24_, 
        nextA_20__23_, nextA_20__22_, nextA_20__21_, nextA_20__20_, 
        nextA_20__19_, nextA_20__18_, nextA_20__17_, nextA_20__16_, 
        nextA_20__15_, nextA_20__14_, nextA_20__13_, nextA_20__12_, 
        nextA_20__11_, nextA_20__10_, nextA_20__9_, nextA_20__8_, nextA_20__7_, 
        nextA_20__6_, nextA_20__5_, nextA_20__4_, nextA_20__3_, nextA_20__2_, 
        nextA_20__1_, nextA_20__0_}), .nextQ({nextQ_20__31_, nextQ_20__30_, 
        nextQ_20__29_, nextQ_20__28_, nextQ_20__27_, nextQ_20__26_, 
        nextQ_20__25_, nextQ_20__24_, nextQ_20__23_, nextQ_20__22_, 
        nextQ_20__21_, nextQ_20__20_, nextQ_20__19_, nextQ_20__18_, 
        nextQ_20__17_, nextQ_20__16_, nextQ_20__15_, nextQ_20__14_, 
        nextQ_20__13_, nextQ_20__12_, nextQ_20__11_, nextQ_20__10_, 
        nextQ_20__9_, nextQ_20__8_, nextQ_20__7_, nextQ_20__6_, nextQ_20__5_, 
        nextQ_20__4_, nextQ_20__3_, nextQ_20__2_, nextQ_20__1_, nextQ_20__0_}), 
        .nextQ_1(q_1[20]) );
  BoothStep_12 booth_instances_20__stepX ( .a({nextA_20__31_, nextA_20__30_, 
        nextA_20__29_, nextA_20__28_, nextA_20__27_, nextA_20__26_, 
        nextA_20__25_, nextA_20__24_, nextA_20__23_, nextA_20__22_, 
        nextA_20__21_, nextA_20__20_, nextA_20__19_, nextA_20__18_, 
        nextA_20__17_, nextA_20__16_, nextA_20__15_, nextA_20__14_, 
        nextA_20__13_, nextA_20__12_, nextA_20__11_, nextA_20__10_, 
        nextA_20__9_, nextA_20__8_, nextA_20__7_, nextA_20__6_, nextA_20__5_, 
        nextA_20__4_, nextA_20__3_, nextA_20__2_, nextA_20__1_, nextA_20__0_}), 
        .q({nextQ_20__31_, nextQ_20__30_, nextQ_20__29_, nextQ_20__28_, 
        nextQ_20__27_, nextQ_20__26_, nextQ_20__25_, nextQ_20__24_, 
        nextQ_20__23_, nextQ_20__22_, nextQ_20__21_, nextQ_20__20_, 
        nextQ_20__19_, nextQ_20__18_, nextQ_20__17_, nextQ_20__16_, 
        nextQ_20__15_, nextQ_20__14_, nextQ_20__13_, nextQ_20__12_, 
        nextQ_20__11_, nextQ_20__10_, nextQ_20__9_, nextQ_20__8_, nextQ_20__7_, 
        nextQ_20__6_, nextQ_20__5_, nextQ_20__4_, nextQ_20__3_, nextQ_20__2_, 
        nextQ_20__1_, nextQ_20__0_}), .m(a), .q_1(q_1[20]), .nextA({
        nextA_21__31_, nextA_21__30_, nextA_21__29_, nextA_21__28_, 
        nextA_21__27_, nextA_21__26_, nextA_21__25_, nextA_21__24_, 
        nextA_21__23_, nextA_21__22_, nextA_21__21_, nextA_21__20_, 
        nextA_21__19_, nextA_21__18_, nextA_21__17_, nextA_21__16_, 
        nextA_21__15_, nextA_21__14_, nextA_21__13_, nextA_21__12_, 
        nextA_21__11_, nextA_21__10_, nextA_21__9_, nextA_21__8_, nextA_21__7_, 
        nextA_21__6_, nextA_21__5_, nextA_21__4_, nextA_21__3_, nextA_21__2_, 
        nextA_21__1_, nextA_21__0_}), .nextQ({nextQ_21__31_, nextQ_21__30_, 
        nextQ_21__29_, nextQ_21__28_, nextQ_21__27_, nextQ_21__26_, 
        nextQ_21__25_, nextQ_21__24_, nextQ_21__23_, nextQ_21__22_, 
        nextQ_21__21_, nextQ_21__20_, nextQ_21__19_, nextQ_21__18_, 
        nextQ_21__17_, nextQ_21__16_, nextQ_21__15_, nextQ_21__14_, 
        nextQ_21__13_, nextQ_21__12_, nextQ_21__11_, nextQ_21__10_, 
        nextQ_21__9_, nextQ_21__8_, nextQ_21__7_, nextQ_21__6_, nextQ_21__5_, 
        nextQ_21__4_, nextQ_21__3_, nextQ_21__2_, nextQ_21__1_, nextQ_21__0_}), 
        .nextQ_1(q_1[21]) );
  BoothStep_11 booth_instances_21__stepX ( .a({nextA_21__31_, nextA_21__30_, 
        nextA_21__29_, nextA_21__28_, nextA_21__27_, nextA_21__26_, 
        nextA_21__25_, nextA_21__24_, nextA_21__23_, nextA_21__22_, 
        nextA_21__21_, nextA_21__20_, nextA_21__19_, nextA_21__18_, 
        nextA_21__17_, nextA_21__16_, nextA_21__15_, nextA_21__14_, 
        nextA_21__13_, nextA_21__12_, nextA_21__11_, nextA_21__10_, 
        nextA_21__9_, nextA_21__8_, nextA_21__7_, nextA_21__6_, nextA_21__5_, 
        nextA_21__4_, nextA_21__3_, nextA_21__2_, nextA_21__1_, nextA_21__0_}), 
        .q({nextQ_21__31_, nextQ_21__30_, nextQ_21__29_, nextQ_21__28_, 
        nextQ_21__27_, nextQ_21__26_, nextQ_21__25_, nextQ_21__24_, 
        nextQ_21__23_, nextQ_21__22_, nextQ_21__21_, nextQ_21__20_, 
        nextQ_21__19_, nextQ_21__18_, nextQ_21__17_, nextQ_21__16_, 
        nextQ_21__15_, nextQ_21__14_, nextQ_21__13_, nextQ_21__12_, 
        nextQ_21__11_, nextQ_21__10_, nextQ_21__9_, nextQ_21__8_, nextQ_21__7_, 
        nextQ_21__6_, nextQ_21__5_, nextQ_21__4_, nextQ_21__3_, nextQ_21__2_, 
        nextQ_21__1_, nextQ_21__0_}), .m(a), .q_1(q_1[21]), .nextA({
        nextA_22__31_, nextA_22__30_, nextA_22__29_, nextA_22__28_, 
        nextA_22__27_, nextA_22__26_, nextA_22__25_, nextA_22__24_, 
        nextA_22__23_, nextA_22__22_, nextA_22__21_, nextA_22__20_, 
        nextA_22__19_, nextA_22__18_, nextA_22__17_, nextA_22__16_, 
        nextA_22__15_, nextA_22__14_, nextA_22__13_, nextA_22__12_, 
        nextA_22__11_, nextA_22__10_, nextA_22__9_, nextA_22__8_, nextA_22__7_, 
        nextA_22__6_, nextA_22__5_, nextA_22__4_, nextA_22__3_, nextA_22__2_, 
        nextA_22__1_, nextA_22__0_}), .nextQ({nextQ_22__31_, nextQ_22__30_, 
        nextQ_22__29_, nextQ_22__28_, nextQ_22__27_, nextQ_22__26_, 
        nextQ_22__25_, nextQ_22__24_, nextQ_22__23_, nextQ_22__22_, 
        nextQ_22__21_, nextQ_22__20_, nextQ_22__19_, nextQ_22__18_, 
        nextQ_22__17_, nextQ_22__16_, nextQ_22__15_, nextQ_22__14_, 
        nextQ_22__13_, nextQ_22__12_, nextQ_22__11_, nextQ_22__10_, 
        nextQ_22__9_, nextQ_22__8_, nextQ_22__7_, nextQ_22__6_, nextQ_22__5_, 
        nextQ_22__4_, nextQ_22__3_, nextQ_22__2_, nextQ_22__1_, nextQ_22__0_}), 
        .nextQ_1(q_1[22]) );
  BoothStep_10 booth_instances_22__stepX ( .a({nextA_22__31_, nextA_22__30_, 
        nextA_22__29_, nextA_22__28_, nextA_22__27_, nextA_22__26_, 
        nextA_22__25_, nextA_22__24_, nextA_22__23_, nextA_22__22_, 
        nextA_22__21_, nextA_22__20_, nextA_22__19_, nextA_22__18_, 
        nextA_22__17_, nextA_22__16_, nextA_22__15_, nextA_22__14_, 
        nextA_22__13_, nextA_22__12_, nextA_22__11_, nextA_22__10_, 
        nextA_22__9_, nextA_22__8_, nextA_22__7_, nextA_22__6_, nextA_22__5_, 
        nextA_22__4_, nextA_22__3_, nextA_22__2_, nextA_22__1_, nextA_22__0_}), 
        .q({nextQ_22__31_, nextQ_22__30_, nextQ_22__29_, nextQ_22__28_, 
        nextQ_22__27_, nextQ_22__26_, nextQ_22__25_, nextQ_22__24_, 
        nextQ_22__23_, nextQ_22__22_, nextQ_22__21_, nextQ_22__20_, 
        nextQ_22__19_, nextQ_22__18_, nextQ_22__17_, nextQ_22__16_, 
        nextQ_22__15_, nextQ_22__14_, nextQ_22__13_, nextQ_22__12_, 
        nextQ_22__11_, nextQ_22__10_, nextQ_22__9_, nextQ_22__8_, nextQ_22__7_, 
        nextQ_22__6_, nextQ_22__5_, nextQ_22__4_, nextQ_22__3_, nextQ_22__2_, 
        nextQ_22__1_, nextQ_22__0_}), .m(a), .q_1(q_1[22]), .nextA({
        nextA_23__31_, nextA_23__30_, nextA_23__29_, nextA_23__28_, 
        nextA_23__27_, nextA_23__26_, nextA_23__25_, nextA_23__24_, 
        nextA_23__23_, nextA_23__22_, nextA_23__21_, nextA_23__20_, 
        nextA_23__19_, nextA_23__18_, nextA_23__17_, nextA_23__16_, 
        nextA_23__15_, nextA_23__14_, nextA_23__13_, nextA_23__12_, 
        nextA_23__11_, nextA_23__10_, nextA_23__9_, nextA_23__8_, nextA_23__7_, 
        nextA_23__6_, nextA_23__5_, nextA_23__4_, nextA_23__3_, nextA_23__2_, 
        nextA_23__1_, nextA_23__0_}), .nextQ({nextQ_23__31_, nextQ_23__30_, 
        nextQ_23__29_, nextQ_23__28_, nextQ_23__27_, nextQ_23__26_, 
        nextQ_23__25_, nextQ_23__24_, nextQ_23__23_, nextQ_23__22_, 
        nextQ_23__21_, nextQ_23__20_, nextQ_23__19_, nextQ_23__18_, 
        nextQ_23__17_, nextQ_23__16_, nextQ_23__15_, nextQ_23__14_, 
        nextQ_23__13_, nextQ_23__12_, nextQ_23__11_, nextQ_23__10_, 
        nextQ_23__9_, nextQ_23__8_, nextQ_23__7_, nextQ_23__6_, nextQ_23__5_, 
        nextQ_23__4_, nextQ_23__3_, nextQ_23__2_, nextQ_23__1_, nextQ_23__0_}), 
        .nextQ_1(q_1[23]) );
  BoothStep_9 booth_instances_23__stepX ( .a({nextA_23__31_, nextA_23__30_, 
        nextA_23__29_, nextA_23__28_, nextA_23__27_, nextA_23__26_, 
        nextA_23__25_, nextA_23__24_, nextA_23__23_, nextA_23__22_, 
        nextA_23__21_, nextA_23__20_, nextA_23__19_, nextA_23__18_, 
        nextA_23__17_, nextA_23__16_, nextA_23__15_, nextA_23__14_, 
        nextA_23__13_, nextA_23__12_, nextA_23__11_, nextA_23__10_, 
        nextA_23__9_, nextA_23__8_, nextA_23__7_, nextA_23__6_, nextA_23__5_, 
        nextA_23__4_, nextA_23__3_, nextA_23__2_, nextA_23__1_, nextA_23__0_}), 
        .q({nextQ_23__31_, nextQ_23__30_, nextQ_23__29_, nextQ_23__28_, 
        nextQ_23__27_, nextQ_23__26_, nextQ_23__25_, nextQ_23__24_, 
        nextQ_23__23_, nextQ_23__22_, nextQ_23__21_, nextQ_23__20_, 
        nextQ_23__19_, nextQ_23__18_, nextQ_23__17_, nextQ_23__16_, 
        nextQ_23__15_, nextQ_23__14_, nextQ_23__13_, nextQ_23__12_, 
        nextQ_23__11_, nextQ_23__10_, nextQ_23__9_, nextQ_23__8_, nextQ_23__7_, 
        nextQ_23__6_, nextQ_23__5_, nextQ_23__4_, nextQ_23__3_, nextQ_23__2_, 
        nextQ_23__1_, nextQ_23__0_}), .m(a), .q_1(q_1[23]), .nextA({
        nextA_24__31_, nextA_24__30_, nextA_24__29_, nextA_24__28_, 
        nextA_24__27_, nextA_24__26_, nextA_24__25_, nextA_24__24_, 
        nextA_24__23_, nextA_24__22_, nextA_24__21_, nextA_24__20_, 
        nextA_24__19_, nextA_24__18_, nextA_24__17_, nextA_24__16_, 
        nextA_24__15_, nextA_24__14_, nextA_24__13_, nextA_24__12_, 
        nextA_24__11_, nextA_24__10_, nextA_24__9_, nextA_24__8_, nextA_24__7_, 
        nextA_24__6_, nextA_24__5_, nextA_24__4_, nextA_24__3_, nextA_24__2_, 
        nextA_24__1_, nextA_24__0_}), .nextQ({nextQ_24__31_, nextQ_24__30_, 
        nextQ_24__29_, nextQ_24__28_, nextQ_24__27_, nextQ_24__26_, 
        nextQ_24__25_, nextQ_24__24_, nextQ_24__23_, nextQ_24__22_, 
        nextQ_24__21_, nextQ_24__20_, nextQ_24__19_, nextQ_24__18_, 
        nextQ_24__17_, nextQ_24__16_, nextQ_24__15_, nextQ_24__14_, 
        nextQ_24__13_, nextQ_24__12_, nextQ_24__11_, nextQ_24__10_, 
        nextQ_24__9_, nextQ_24__8_, nextQ_24__7_, nextQ_24__6_, nextQ_24__5_, 
        nextQ_24__4_, nextQ_24__3_, nextQ_24__2_, nextQ_24__1_, nextQ_24__0_}), 
        .nextQ_1(q_1[24]) );
  BoothStep_8 booth_instances_24__stepX ( .a({nextA_24__31_, nextA_24__30_, 
        nextA_24__29_, nextA_24__28_, nextA_24__27_, nextA_24__26_, 
        nextA_24__25_, nextA_24__24_, nextA_24__23_, nextA_24__22_, 
        nextA_24__21_, nextA_24__20_, nextA_24__19_, nextA_24__18_, 
        nextA_24__17_, nextA_24__16_, nextA_24__15_, nextA_24__14_, 
        nextA_24__13_, nextA_24__12_, nextA_24__11_, nextA_24__10_, 
        nextA_24__9_, nextA_24__8_, nextA_24__7_, nextA_24__6_, nextA_24__5_, 
        nextA_24__4_, nextA_24__3_, nextA_24__2_, nextA_24__1_, nextA_24__0_}), 
        .q({nextQ_24__31_, nextQ_24__30_, nextQ_24__29_, nextQ_24__28_, 
        nextQ_24__27_, nextQ_24__26_, nextQ_24__25_, nextQ_24__24_, 
        nextQ_24__23_, nextQ_24__22_, nextQ_24__21_, nextQ_24__20_, 
        nextQ_24__19_, nextQ_24__18_, nextQ_24__17_, nextQ_24__16_, 
        nextQ_24__15_, nextQ_24__14_, nextQ_24__13_, nextQ_24__12_, 
        nextQ_24__11_, nextQ_24__10_, nextQ_24__9_, nextQ_24__8_, nextQ_24__7_, 
        nextQ_24__6_, nextQ_24__5_, nextQ_24__4_, nextQ_24__3_, nextQ_24__2_, 
        nextQ_24__1_, nextQ_24__0_}), .m(a), .q_1(q_1[24]), .nextA({
        nextA_25__31_, nextA_25__30_, nextA_25__29_, nextA_25__28_, 
        nextA_25__27_, nextA_25__26_, nextA_25__25_, nextA_25__24_, 
        nextA_25__23_, nextA_25__22_, nextA_25__21_, nextA_25__20_, 
        nextA_25__19_, nextA_25__18_, nextA_25__17_, nextA_25__16_, 
        nextA_25__15_, nextA_25__14_, nextA_25__13_, nextA_25__12_, 
        nextA_25__11_, nextA_25__10_, nextA_25__9_, nextA_25__8_, nextA_25__7_, 
        nextA_25__6_, nextA_25__5_, nextA_25__4_, nextA_25__3_, nextA_25__2_, 
        nextA_25__1_, nextA_25__0_}), .nextQ({nextQ_25__31_, nextQ_25__30_, 
        nextQ_25__29_, nextQ_25__28_, nextQ_25__27_, nextQ_25__26_, 
        nextQ_25__25_, nextQ_25__24_, nextQ_25__23_, nextQ_25__22_, 
        nextQ_25__21_, nextQ_25__20_, nextQ_25__19_, nextQ_25__18_, 
        nextQ_25__17_, nextQ_25__16_, nextQ_25__15_, nextQ_25__14_, 
        nextQ_25__13_, nextQ_25__12_, nextQ_25__11_, nextQ_25__10_, 
        nextQ_25__9_, nextQ_25__8_, nextQ_25__7_, nextQ_25__6_, nextQ_25__5_, 
        nextQ_25__4_, nextQ_25__3_, nextQ_25__2_, nextQ_25__1_, nextQ_25__0_}), 
        .nextQ_1(q_1[25]) );
  BoothStep_7 booth_instances_25__stepX ( .a({nextA_25__31_, nextA_25__30_, 
        nextA_25__29_, nextA_25__28_, nextA_25__27_, nextA_25__26_, 
        nextA_25__25_, nextA_25__24_, nextA_25__23_, nextA_25__22_, 
        nextA_25__21_, nextA_25__20_, nextA_25__19_, nextA_25__18_, 
        nextA_25__17_, nextA_25__16_, nextA_25__15_, nextA_25__14_, 
        nextA_25__13_, nextA_25__12_, nextA_25__11_, nextA_25__10_, 
        nextA_25__9_, nextA_25__8_, nextA_25__7_, nextA_25__6_, nextA_25__5_, 
        nextA_25__4_, nextA_25__3_, nextA_25__2_, nextA_25__1_, nextA_25__0_}), 
        .q({nextQ_25__31_, nextQ_25__30_, nextQ_25__29_, nextQ_25__28_, 
        nextQ_25__27_, nextQ_25__26_, nextQ_25__25_, nextQ_25__24_, 
        nextQ_25__23_, nextQ_25__22_, nextQ_25__21_, nextQ_25__20_, 
        nextQ_25__19_, nextQ_25__18_, nextQ_25__17_, nextQ_25__16_, 
        nextQ_25__15_, nextQ_25__14_, nextQ_25__13_, nextQ_25__12_, 
        nextQ_25__11_, nextQ_25__10_, nextQ_25__9_, nextQ_25__8_, nextQ_25__7_, 
        nextQ_25__6_, nextQ_25__5_, nextQ_25__4_, nextQ_25__3_, nextQ_25__2_, 
        nextQ_25__1_, nextQ_25__0_}), .m(a), .q_1(q_1[25]), .nextA({
        nextA_26__31_, nextA_26__30_, nextA_26__29_, nextA_26__28_, 
        nextA_26__27_, nextA_26__26_, nextA_26__25_, nextA_26__24_, 
        nextA_26__23_, nextA_26__22_, nextA_26__21_, nextA_26__20_, 
        nextA_26__19_, nextA_26__18_, nextA_26__17_, nextA_26__16_, 
        nextA_26__15_, nextA_26__14_, nextA_26__13_, nextA_26__12_, 
        nextA_26__11_, nextA_26__10_, nextA_26__9_, nextA_26__8_, nextA_26__7_, 
        nextA_26__6_, nextA_26__5_, nextA_26__4_, nextA_26__3_, nextA_26__2_, 
        nextA_26__1_, nextA_26__0_}), .nextQ({nextQ_26__31_, nextQ_26__30_, 
        nextQ_26__29_, nextQ_26__28_, nextQ_26__27_, nextQ_26__26_, 
        nextQ_26__25_, nextQ_26__24_, nextQ_26__23_, nextQ_26__22_, 
        nextQ_26__21_, nextQ_26__20_, nextQ_26__19_, nextQ_26__18_, 
        nextQ_26__17_, nextQ_26__16_, nextQ_26__15_, nextQ_26__14_, 
        nextQ_26__13_, nextQ_26__12_, nextQ_26__11_, nextQ_26__10_, 
        nextQ_26__9_, nextQ_26__8_, nextQ_26__7_, nextQ_26__6_, nextQ_26__5_, 
        nextQ_26__4_, nextQ_26__3_, nextQ_26__2_, nextQ_26__1_, nextQ_26__0_}), 
        .nextQ_1(q_1[26]) );
  BoothStep_6 booth_instances_26__stepX ( .a({nextA_26__31_, nextA_26__30_, 
        nextA_26__29_, nextA_26__28_, nextA_26__27_, nextA_26__26_, 
        nextA_26__25_, nextA_26__24_, nextA_26__23_, nextA_26__22_, 
        nextA_26__21_, nextA_26__20_, nextA_26__19_, nextA_26__18_, 
        nextA_26__17_, nextA_26__16_, nextA_26__15_, nextA_26__14_, 
        nextA_26__13_, nextA_26__12_, nextA_26__11_, nextA_26__10_, 
        nextA_26__9_, nextA_26__8_, nextA_26__7_, nextA_26__6_, nextA_26__5_, 
        nextA_26__4_, nextA_26__3_, nextA_26__2_, nextA_26__1_, nextA_26__0_}), 
        .q({nextQ_26__31_, nextQ_26__30_, nextQ_26__29_, nextQ_26__28_, 
        nextQ_26__27_, nextQ_26__26_, nextQ_26__25_, nextQ_26__24_, 
        nextQ_26__23_, nextQ_26__22_, nextQ_26__21_, nextQ_26__20_, 
        nextQ_26__19_, nextQ_26__18_, nextQ_26__17_, nextQ_26__16_, 
        nextQ_26__15_, nextQ_26__14_, nextQ_26__13_, nextQ_26__12_, 
        nextQ_26__11_, nextQ_26__10_, nextQ_26__9_, nextQ_26__8_, nextQ_26__7_, 
        nextQ_26__6_, nextQ_26__5_, nextQ_26__4_, nextQ_26__3_, nextQ_26__2_, 
        nextQ_26__1_, nextQ_26__0_}), .m(a), .q_1(q_1[26]), .nextA({
        nextA_27__31_, nextA_27__30_, nextA_27__29_, nextA_27__28_, 
        nextA_27__27_, nextA_27__26_, nextA_27__25_, nextA_27__24_, 
        nextA_27__23_, nextA_27__22_, nextA_27__21_, nextA_27__20_, 
        nextA_27__19_, nextA_27__18_, nextA_27__17_, nextA_27__16_, 
        nextA_27__15_, nextA_27__14_, nextA_27__13_, nextA_27__12_, 
        nextA_27__11_, nextA_27__10_, nextA_27__9_, nextA_27__8_, nextA_27__7_, 
        nextA_27__6_, nextA_27__5_, nextA_27__4_, nextA_27__3_, nextA_27__2_, 
        nextA_27__1_, nextA_27__0_}), .nextQ({nextQ_27__31_, nextQ_27__30_, 
        nextQ_27__29_, nextQ_27__28_, nextQ_27__27_, nextQ_27__26_, 
        nextQ_27__25_, nextQ_27__24_, nextQ_27__23_, nextQ_27__22_, 
        nextQ_27__21_, nextQ_27__20_, nextQ_27__19_, nextQ_27__18_, 
        nextQ_27__17_, nextQ_27__16_, nextQ_27__15_, nextQ_27__14_, 
        nextQ_27__13_, nextQ_27__12_, nextQ_27__11_, nextQ_27__10_, 
        nextQ_27__9_, nextQ_27__8_, nextQ_27__7_, nextQ_27__6_, nextQ_27__5_, 
        nextQ_27__4_, nextQ_27__3_, nextQ_27__2_, nextQ_27__1_, nextQ_27__0_}), 
        .nextQ_1(q_1[27]) );
  BoothStep_5 booth_instances_27__stepX ( .a({nextA_27__31_, nextA_27__30_, 
        nextA_27__29_, nextA_27__28_, nextA_27__27_, nextA_27__26_, 
        nextA_27__25_, nextA_27__24_, nextA_27__23_, nextA_27__22_, 
        nextA_27__21_, nextA_27__20_, nextA_27__19_, nextA_27__18_, 
        nextA_27__17_, nextA_27__16_, nextA_27__15_, nextA_27__14_, 
        nextA_27__13_, nextA_27__12_, nextA_27__11_, nextA_27__10_, 
        nextA_27__9_, nextA_27__8_, nextA_27__7_, nextA_27__6_, nextA_27__5_, 
        nextA_27__4_, nextA_27__3_, nextA_27__2_, nextA_27__1_, nextA_27__0_}), 
        .q({nextQ_27__31_, nextQ_27__30_, nextQ_27__29_, nextQ_27__28_, 
        nextQ_27__27_, nextQ_27__26_, nextQ_27__25_, nextQ_27__24_, 
        nextQ_27__23_, nextQ_27__22_, nextQ_27__21_, nextQ_27__20_, 
        nextQ_27__19_, nextQ_27__18_, nextQ_27__17_, nextQ_27__16_, 
        nextQ_27__15_, nextQ_27__14_, nextQ_27__13_, nextQ_27__12_, 
        nextQ_27__11_, nextQ_27__10_, nextQ_27__9_, nextQ_27__8_, nextQ_27__7_, 
        nextQ_27__6_, nextQ_27__5_, nextQ_27__4_, nextQ_27__3_, nextQ_27__2_, 
        nextQ_27__1_, nextQ_27__0_}), .m(a), .q_1(q_1[27]), .nextA({
        nextA_28__31_, nextA_28__30_, nextA_28__29_, nextA_28__28_, 
        nextA_28__27_, nextA_28__26_, nextA_28__25_, nextA_28__24_, 
        nextA_28__23_, nextA_28__22_, nextA_28__21_, nextA_28__20_, 
        nextA_28__19_, nextA_28__18_, nextA_28__17_, nextA_28__16_, 
        nextA_28__15_, nextA_28__14_, nextA_28__13_, nextA_28__12_, 
        nextA_28__11_, nextA_28__10_, nextA_28__9_, nextA_28__8_, nextA_28__7_, 
        nextA_28__6_, nextA_28__5_, nextA_28__4_, nextA_28__3_, nextA_28__2_, 
        nextA_28__1_, nextA_28__0_}), .nextQ({nextQ_28__31_, nextQ_28__30_, 
        nextQ_28__29_, nextQ_28__28_, nextQ_28__27_, nextQ_28__26_, 
        nextQ_28__25_, nextQ_28__24_, nextQ_28__23_, nextQ_28__22_, 
        nextQ_28__21_, nextQ_28__20_, nextQ_28__19_, nextQ_28__18_, 
        nextQ_28__17_, nextQ_28__16_, nextQ_28__15_, nextQ_28__14_, 
        nextQ_28__13_, nextQ_28__12_, nextQ_28__11_, nextQ_28__10_, 
        nextQ_28__9_, nextQ_28__8_, nextQ_28__7_, nextQ_28__6_, nextQ_28__5_, 
        nextQ_28__4_, nextQ_28__3_, nextQ_28__2_, nextQ_28__1_, nextQ_28__0_}), 
        .nextQ_1(q_1[28]) );
  BoothStep_4 booth_instances_28__stepX ( .a({nextA_28__31_, nextA_28__30_, 
        nextA_28__29_, nextA_28__28_, nextA_28__27_, nextA_28__26_, 
        nextA_28__25_, nextA_28__24_, nextA_28__23_, nextA_28__22_, 
        nextA_28__21_, nextA_28__20_, nextA_28__19_, nextA_28__18_, 
        nextA_28__17_, nextA_28__16_, nextA_28__15_, nextA_28__14_, 
        nextA_28__13_, nextA_28__12_, nextA_28__11_, nextA_28__10_, 
        nextA_28__9_, nextA_28__8_, nextA_28__7_, nextA_28__6_, nextA_28__5_, 
        nextA_28__4_, nextA_28__3_, nextA_28__2_, nextA_28__1_, nextA_28__0_}), 
        .q({nextQ_28__31_, nextQ_28__30_, nextQ_28__29_, nextQ_28__28_, 
        nextQ_28__27_, nextQ_28__26_, nextQ_28__25_, nextQ_28__24_, 
        nextQ_28__23_, nextQ_28__22_, nextQ_28__21_, nextQ_28__20_, 
        nextQ_28__19_, nextQ_28__18_, nextQ_28__17_, nextQ_28__16_, 
        nextQ_28__15_, nextQ_28__14_, nextQ_28__13_, nextQ_28__12_, 
        nextQ_28__11_, nextQ_28__10_, nextQ_28__9_, nextQ_28__8_, nextQ_28__7_, 
        nextQ_28__6_, nextQ_28__5_, nextQ_28__4_, nextQ_28__3_, nextQ_28__2_, 
        nextQ_28__1_, nextQ_28__0_}), .m(a), .q_1(q_1[28]), .nextA({
        nextA_29__31_, nextA_29__30_, nextA_29__29_, nextA_29__28_, 
        nextA_29__27_, nextA_29__26_, nextA_29__25_, nextA_29__24_, 
        nextA_29__23_, nextA_29__22_, nextA_29__21_, nextA_29__20_, 
        nextA_29__19_, nextA_29__18_, nextA_29__17_, nextA_29__16_, 
        nextA_29__15_, nextA_29__14_, nextA_29__13_, nextA_29__12_, 
        nextA_29__11_, nextA_29__10_, nextA_29__9_, nextA_29__8_, nextA_29__7_, 
        nextA_29__6_, nextA_29__5_, nextA_29__4_, nextA_29__3_, nextA_29__2_, 
        nextA_29__1_, nextA_29__0_}), .nextQ({nextQ_29__31_, nextQ_29__30_, 
        nextQ_29__29_, nextQ_29__28_, nextQ_29__27_, nextQ_29__26_, 
        nextQ_29__25_, nextQ_29__24_, nextQ_29__23_, nextQ_29__22_, 
        nextQ_29__21_, nextQ_29__20_, nextQ_29__19_, nextQ_29__18_, 
        nextQ_29__17_, nextQ_29__16_, nextQ_29__15_, nextQ_29__14_, 
        nextQ_29__13_, nextQ_29__12_, nextQ_29__11_, nextQ_29__10_, 
        nextQ_29__9_, nextQ_29__8_, nextQ_29__7_, nextQ_29__6_, nextQ_29__5_, 
        nextQ_29__4_, nextQ_29__3_, nextQ_29__2_, nextQ_29__1_, nextQ_29__0_}), 
        .nextQ_1(q_1[29]) );
  BoothStep_3 booth_instances_29__stepX ( .a({nextA_29__31_, nextA_29__30_, 
        nextA_29__29_, nextA_29__28_, nextA_29__27_, nextA_29__26_, 
        nextA_29__25_, nextA_29__24_, nextA_29__23_, nextA_29__22_, 
        nextA_29__21_, nextA_29__20_, nextA_29__19_, nextA_29__18_, 
        nextA_29__17_, nextA_29__16_, nextA_29__15_, nextA_29__14_, 
        nextA_29__13_, nextA_29__12_, nextA_29__11_, nextA_29__10_, 
        nextA_29__9_, nextA_29__8_, nextA_29__7_, nextA_29__6_, nextA_29__5_, 
        nextA_29__4_, nextA_29__3_, nextA_29__2_, nextA_29__1_, nextA_29__0_}), 
        .q({nextQ_29__31_, nextQ_29__30_, nextQ_29__29_, nextQ_29__28_, 
        nextQ_29__27_, nextQ_29__26_, nextQ_29__25_, nextQ_29__24_, 
        nextQ_29__23_, nextQ_29__22_, nextQ_29__21_, nextQ_29__20_, 
        nextQ_29__19_, nextQ_29__18_, nextQ_29__17_, nextQ_29__16_, 
        nextQ_29__15_, nextQ_29__14_, nextQ_29__13_, nextQ_29__12_, 
        nextQ_29__11_, nextQ_29__10_, nextQ_29__9_, nextQ_29__8_, nextQ_29__7_, 
        nextQ_29__6_, nextQ_29__5_, nextQ_29__4_, nextQ_29__3_, nextQ_29__2_, 
        nextQ_29__1_, nextQ_29__0_}), .m(a), .q_1(q_1[29]), .nextA({
        nextA_30__31_, nextA_30__30_, nextA_30__29_, nextA_30__28_, 
        nextA_30__27_, nextA_30__26_, nextA_30__25_, nextA_30__24_, 
        nextA_30__23_, nextA_30__22_, nextA_30__21_, nextA_30__20_, 
        nextA_30__19_, nextA_30__18_, nextA_30__17_, nextA_30__16_, 
        nextA_30__15_, nextA_30__14_, nextA_30__13_, nextA_30__12_, 
        nextA_30__11_, nextA_30__10_, nextA_30__9_, nextA_30__8_, nextA_30__7_, 
        nextA_30__6_, nextA_30__5_, nextA_30__4_, nextA_30__3_, nextA_30__2_, 
        nextA_30__1_, nextA_30__0_}), .nextQ({nextQ_30__31_, nextQ_30__30_, 
        nextQ_30__29_, nextQ_30__28_, nextQ_30__27_, nextQ_30__26_, 
        nextQ_30__25_, nextQ_30__24_, nextQ_30__23_, nextQ_30__22_, 
        nextQ_30__21_, nextQ_30__20_, nextQ_30__19_, nextQ_30__18_, 
        nextQ_30__17_, nextQ_30__16_, nextQ_30__15_, nextQ_30__14_, 
        nextQ_30__13_, nextQ_30__12_, nextQ_30__11_, nextQ_30__10_, 
        nextQ_30__9_, nextQ_30__8_, nextQ_30__7_, nextQ_30__6_, nextQ_30__5_, 
        nextQ_30__4_, nextQ_30__3_, nextQ_30__2_, nextQ_30__1_, nextQ_30__0_}), 
        .nextQ_1(q_1[30]) );
  BoothStep_2 booth_instances_30__stepX ( .a({nextA_30__31_, nextA_30__30_, 
        nextA_30__29_, nextA_30__28_, nextA_30__27_, nextA_30__26_, 
        nextA_30__25_, nextA_30__24_, nextA_30__23_, nextA_30__22_, 
        nextA_30__21_, nextA_30__20_, nextA_30__19_, nextA_30__18_, 
        nextA_30__17_, nextA_30__16_, nextA_30__15_, nextA_30__14_, 
        nextA_30__13_, nextA_30__12_, nextA_30__11_, nextA_30__10_, 
        nextA_30__9_, nextA_30__8_, nextA_30__7_, nextA_30__6_, nextA_30__5_, 
        nextA_30__4_, nextA_30__3_, nextA_30__2_, nextA_30__1_, nextA_30__0_}), 
        .q({nextQ_30__31_, nextQ_30__30_, nextQ_30__29_, nextQ_30__28_, 
        nextQ_30__27_, nextQ_30__26_, nextQ_30__25_, nextQ_30__24_, 
        nextQ_30__23_, nextQ_30__22_, nextQ_30__21_, nextQ_30__20_, 
        nextQ_30__19_, nextQ_30__18_, nextQ_30__17_, nextQ_30__16_, 
        nextQ_30__15_, nextQ_30__14_, nextQ_30__13_, nextQ_30__12_, 
        nextQ_30__11_, nextQ_30__10_, nextQ_30__9_, nextQ_30__8_, nextQ_30__7_, 
        nextQ_30__6_, nextQ_30__5_, nextQ_30__4_, nextQ_30__3_, nextQ_30__2_, 
        nextQ_30__1_, nextQ_30__0_}), .m(a), .q_1(q_1[30]), .nextA({
        nextA_31__31_, nextA_31__30_, nextA_31__29_, nextA_31__28_, 
        nextA_31__27_, nextA_31__26_, nextA_31__25_, nextA_31__24_, 
        nextA_31__23_, nextA_31__22_, nextA_31__21_, nextA_31__20_, 
        nextA_31__19_, nextA_31__18_, nextA_31__17_, nextA_31__16_, 
        nextA_31__15_, nextA_31__14_, nextA_31__13_, nextA_31__12_, 
        nextA_31__11_, nextA_31__10_, nextA_31__9_, nextA_31__8_, nextA_31__7_, 
        nextA_31__6_, nextA_31__5_, nextA_31__4_, nextA_31__3_, nextA_31__2_, 
        nextA_31__1_, nextA_31__0_}), .nextQ({nextQ_31__31_, nextQ_31__30_, 
        nextQ_31__29_, nextQ_31__28_, nextQ_31__27_, nextQ_31__26_, 
        nextQ_31__25_, nextQ_31__24_, nextQ_31__23_, nextQ_31__22_, 
        nextQ_31__21_, nextQ_31__20_, nextQ_31__19_, nextQ_31__18_, 
        nextQ_31__17_, nextQ_31__16_, nextQ_31__15_, nextQ_31__14_, 
        nextQ_31__13_, nextQ_31__12_, nextQ_31__11_, nextQ_31__10_, 
        nextQ_31__9_, nextQ_31__8_, nextQ_31__7_, nextQ_31__6_, nextQ_31__5_, 
        nextQ_31__4_, nextQ_31__3_, nextQ_31__2_, nextQ_31__1_, nextQ_31__0_}), 
        .nextQ_1(q_1[31]) );
  BoothStep_1 booth_instances_31__stepX ( .a({nextA_31__31_, nextA_31__30_, 
        nextA_31__29_, nextA_31__28_, nextA_31__27_, nextA_31__26_, 
        nextA_31__25_, nextA_31__24_, nextA_31__23_, nextA_31__22_, 
        nextA_31__21_, nextA_31__20_, nextA_31__19_, nextA_31__18_, 
        nextA_31__17_, nextA_31__16_, nextA_31__15_, nextA_31__14_, 
        nextA_31__13_, nextA_31__12_, nextA_31__11_, nextA_31__10_, 
        nextA_31__9_, nextA_31__8_, nextA_31__7_, nextA_31__6_, nextA_31__5_, 
        nextA_31__4_, nextA_31__3_, nextA_31__2_, nextA_31__1_, nextA_31__0_}), 
        .q({nextQ_31__31_, nextQ_31__30_, nextQ_31__29_, nextQ_31__28_, 
        nextQ_31__27_, nextQ_31__26_, nextQ_31__25_, nextQ_31__24_, 
        nextQ_31__23_, nextQ_31__22_, nextQ_31__21_, nextQ_31__20_, 
        nextQ_31__19_, nextQ_31__18_, nextQ_31__17_, nextQ_31__16_, 
        nextQ_31__15_, nextQ_31__14_, nextQ_31__13_, nextQ_31__12_, 
        nextQ_31__11_, nextQ_31__10_, nextQ_31__9_, nextQ_31__8_, nextQ_31__7_, 
        nextQ_31__6_, nextQ_31__5_, nextQ_31__4_, nextQ_31__3_, nextQ_31__2_, 
        nextQ_31__1_, nextQ_31__0_}), .m(a), .q_1(q_1[31]), .nextA(
        result[63:32]), .nextQ(result[31:0]) );
endmodule


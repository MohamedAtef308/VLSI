
module FullAdder_0 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_33 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_34 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_35 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_36 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_37 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_38 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_39 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_40 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_41 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_42 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_43 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_44 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_45 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_46 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_47 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_48 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_49 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_50 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_51 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_52 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_53 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_54 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_55 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_56 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_57 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_58 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_59 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_60 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_61 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_62 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_63 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_0 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_0 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_63 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_62 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_61 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_60 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_59 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_58 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_57 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_56 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_55 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_54 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_53 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_52 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_51 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_50 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_49 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_48 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_47 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_46 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_45 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_44 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_43 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_42 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_41 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_40 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_39 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_38 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_37 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_36 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_35 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_34 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_33 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), 
        .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module FullAdder_1 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_3 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_4 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_5 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_6 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_7 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_8 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_9 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_10 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_11 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_12 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_13 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_14 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_15 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_16 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_17 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_18 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_19 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_20 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_21 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_22 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_23 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_24 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_25 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_26 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_27 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_28 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_29 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_30 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_31 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_32 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_32_1 ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [30:0] passCout;

  FullAdder_32 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_31 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_30 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_29 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_28 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_27 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_26 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_25 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_24 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_23 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_22 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_21 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_20 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_19 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_18 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_17 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_16 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_15 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_14 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_13 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_12 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_11 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_10 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_9 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_8 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_7 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_6 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_5 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_4 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_3 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_2 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_1 bit63 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), 
        .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[31]), .B(a[31]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[31]), .B(sum[31]), .ZN(n1) );
endmodule


module BoothStep ( a, q, m, q_1, nextA, nextQ, nextQ_1 );
  input [31:0] a;
  input [31:0] q;
  input [31:0] m;
  output [31:0] nextA;
  output [31:0] nextQ;
  input q_1;
  output nextQ_1;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136;
  wire   [31:0] sumAM;
  wire   [31:0] subAM;
  assign nextQ_1 = q[0];
  assign nextQ[30] = q[31];
  assign nextQ[29] = q[30];
  assign nextQ[28] = q[29];
  assign nextQ[27] = q[28];
  assign nextQ[26] = q[27];
  assign nextQ[25] = q[26];
  assign nextQ[24] = q[25];
  assign nextQ[23] = q[24];
  assign nextQ[22] = q[23];
  assign nextQ[21] = q[22];
  assign nextQ[20] = q[21];
  assign nextQ[19] = q[20];
  assign nextQ[18] = q[19];
  assign nextQ[17] = q[18];
  assign nextQ[16] = q[17];
  assign nextQ[15] = q[16];
  assign nextQ[14] = q[15];
  assign nextQ[13] = q[14];
  assign nextQ[12] = q[13];
  assign nextQ[11] = q[12];
  assign nextQ[10] = q[11];
  assign nextQ[9] = q[10];
  assign nextQ[8] = q[9];
  assign nextQ[7] = q[8];
  assign nextQ[6] = q[7];
  assign nextQ[5] = q[6];
  assign nextQ[4] = q[5];
  assign nextQ[3] = q[4];
  assign nextQ[2] = q[3];
  assign nextQ[1] = q[2];
  assign nextQ[0] = q[1];
  assign nextA[31] = nextA[30];

  CRAdder_32_0 sum ( .a(a), .b(m), .cin(1'b0), .sum(sumAM) );
  CRAdder_32_1 sub ( .a(a), .b({n33, n34, n35, n36, n37, n38, n39, n40, n41, 
        n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, 
        n56, n57, n58, n59, n60, n61, n62, n63, n64}), .cin(1'b1), .sum(subAM)
         );
  NOR2_X4 U103 ( .A1(n104), .A2(n102), .ZN(n103) );
  NOR2_X4 U104 ( .A1(n136), .A2(q[0]), .ZN(n102) );
  AND2_X2 U105 ( .A1(q[0]), .A2(n136), .ZN(n104) );
  INV_X1 U106 ( .A(n101), .ZN(nextQ[31]) );
  AOI222_X1 U107 ( .A1(sumAM[0]), .A2(n102), .B1(a[0]), .B2(n103), .C1(
        subAM[0]), .C2(n104), .ZN(n101) );
  INV_X1 U108 ( .A(n105), .ZN(nextA[9]) );
  AOI222_X1 U109 ( .A1(sumAM[10]), .A2(n102), .B1(a[10]), .B2(n103), .C1(
        subAM[10]), .C2(n104), .ZN(n105) );
  INV_X1 U110 ( .A(n106), .ZN(nextA[8]) );
  AOI222_X1 U111 ( .A1(sumAM[9]), .A2(n102), .B1(a[9]), .B2(n103), .C1(
        subAM[9]), .C2(n104), .ZN(n106) );
  INV_X1 U112 ( .A(n107), .ZN(nextA[7]) );
  AOI222_X1 U113 ( .A1(sumAM[8]), .A2(n102), .B1(a[8]), .B2(n103), .C1(
        subAM[8]), .C2(n104), .ZN(n107) );
  INV_X1 U114 ( .A(n108), .ZN(nextA[6]) );
  AOI222_X1 U115 ( .A1(sumAM[7]), .A2(n102), .B1(a[7]), .B2(n103), .C1(
        subAM[7]), .C2(n104), .ZN(n108) );
  INV_X1 U116 ( .A(n109), .ZN(nextA[5]) );
  AOI222_X1 U117 ( .A1(sumAM[6]), .A2(n102), .B1(a[6]), .B2(n103), .C1(
        subAM[6]), .C2(n104), .ZN(n109) );
  INV_X1 U118 ( .A(n110), .ZN(nextA[4]) );
  AOI222_X1 U119 ( .A1(sumAM[5]), .A2(n102), .B1(a[5]), .B2(n103), .C1(
        subAM[5]), .C2(n104), .ZN(n110) );
  INV_X1 U120 ( .A(n111), .ZN(nextA[3]) );
  AOI222_X1 U121 ( .A1(sumAM[4]), .A2(n102), .B1(a[4]), .B2(n103), .C1(
        subAM[4]), .C2(n104), .ZN(n111) );
  INV_X1 U122 ( .A(n112), .ZN(nextA[30]) );
  AOI222_X1 U123 ( .A1(sumAM[31]), .A2(n102), .B1(a[31]), .B2(n103), .C1(
        subAM[31]), .C2(n104), .ZN(n112) );
  INV_X1 U124 ( .A(n113), .ZN(nextA[2]) );
  AOI222_X1 U125 ( .A1(sumAM[3]), .A2(n102), .B1(a[3]), .B2(n103), .C1(
        subAM[3]), .C2(n104), .ZN(n113) );
  INV_X1 U126 ( .A(n114), .ZN(nextA[29]) );
  AOI222_X1 U127 ( .A1(sumAM[30]), .A2(n102), .B1(a[30]), .B2(n103), .C1(
        subAM[30]), .C2(n104), .ZN(n114) );
  INV_X1 U128 ( .A(n115), .ZN(nextA[28]) );
  AOI222_X1 U129 ( .A1(sumAM[29]), .A2(n102), .B1(a[29]), .B2(n103), .C1(
        subAM[29]), .C2(n104), .ZN(n115) );
  INV_X1 U130 ( .A(n116), .ZN(nextA[27]) );
  AOI222_X1 U131 ( .A1(sumAM[28]), .A2(n102), .B1(a[28]), .B2(n103), .C1(
        subAM[28]), .C2(n104), .ZN(n116) );
  INV_X1 U132 ( .A(n117), .ZN(nextA[26]) );
  AOI222_X1 U133 ( .A1(sumAM[27]), .A2(n102), .B1(a[27]), .B2(n103), .C1(
        subAM[27]), .C2(n104), .ZN(n117) );
  INV_X1 U134 ( .A(n118), .ZN(nextA[25]) );
  AOI222_X1 U135 ( .A1(sumAM[26]), .A2(n102), .B1(a[26]), .B2(n103), .C1(
        subAM[26]), .C2(n104), .ZN(n118) );
  INV_X1 U136 ( .A(n119), .ZN(nextA[24]) );
  AOI222_X1 U137 ( .A1(sumAM[25]), .A2(n102), .B1(a[25]), .B2(n103), .C1(
        subAM[25]), .C2(n104), .ZN(n119) );
  INV_X1 U138 ( .A(n120), .ZN(nextA[23]) );
  AOI222_X1 U139 ( .A1(sumAM[24]), .A2(n102), .B1(a[24]), .B2(n103), .C1(
        subAM[24]), .C2(n104), .ZN(n120) );
  INV_X1 U140 ( .A(n121), .ZN(nextA[22]) );
  AOI222_X1 U141 ( .A1(sumAM[23]), .A2(n102), .B1(a[23]), .B2(n103), .C1(
        subAM[23]), .C2(n104), .ZN(n121) );
  INV_X1 U142 ( .A(n122), .ZN(nextA[21]) );
  AOI222_X1 U143 ( .A1(sumAM[22]), .A2(n102), .B1(a[22]), .B2(n103), .C1(
        subAM[22]), .C2(n104), .ZN(n122) );
  INV_X1 U144 ( .A(n123), .ZN(nextA[20]) );
  AOI222_X1 U145 ( .A1(sumAM[21]), .A2(n102), .B1(a[21]), .B2(n103), .C1(
        subAM[21]), .C2(n104), .ZN(n123) );
  INV_X1 U146 ( .A(n124), .ZN(nextA[1]) );
  AOI222_X1 U147 ( .A1(sumAM[2]), .A2(n102), .B1(a[2]), .B2(n103), .C1(
        subAM[2]), .C2(n104), .ZN(n124) );
  INV_X1 U148 ( .A(n125), .ZN(nextA[19]) );
  AOI222_X1 U149 ( .A1(sumAM[20]), .A2(n102), .B1(a[20]), .B2(n103), .C1(
        subAM[20]), .C2(n104), .ZN(n125) );
  INV_X1 U150 ( .A(n126), .ZN(nextA[18]) );
  AOI222_X1 U151 ( .A1(sumAM[19]), .A2(n102), .B1(a[19]), .B2(n103), .C1(
        subAM[19]), .C2(n104), .ZN(n126) );
  INV_X1 U152 ( .A(n127), .ZN(nextA[17]) );
  AOI222_X1 U153 ( .A1(sumAM[18]), .A2(n102), .B1(a[18]), .B2(n103), .C1(
        subAM[18]), .C2(n104), .ZN(n127) );
  INV_X1 U154 ( .A(n128), .ZN(nextA[16]) );
  AOI222_X1 U155 ( .A1(sumAM[17]), .A2(n102), .B1(a[17]), .B2(n103), .C1(
        subAM[17]), .C2(n104), .ZN(n128) );
  INV_X1 U156 ( .A(n129), .ZN(nextA[15]) );
  AOI222_X1 U157 ( .A1(sumAM[16]), .A2(n102), .B1(a[16]), .B2(n103), .C1(
        subAM[16]), .C2(n104), .ZN(n129) );
  INV_X1 U158 ( .A(n130), .ZN(nextA[14]) );
  AOI222_X1 U159 ( .A1(sumAM[15]), .A2(n102), .B1(a[15]), .B2(n103), .C1(
        subAM[15]), .C2(n104), .ZN(n130) );
  INV_X1 U160 ( .A(n131), .ZN(nextA[13]) );
  AOI222_X1 U161 ( .A1(sumAM[14]), .A2(n102), .B1(a[14]), .B2(n103), .C1(
        subAM[14]), .C2(n104), .ZN(n131) );
  INV_X1 U162 ( .A(n132), .ZN(nextA[12]) );
  AOI222_X1 U163 ( .A1(sumAM[13]), .A2(n102), .B1(a[13]), .B2(n103), .C1(
        subAM[13]), .C2(n104), .ZN(n132) );
  INV_X1 U164 ( .A(n133), .ZN(nextA[11]) );
  AOI222_X1 U165 ( .A1(sumAM[12]), .A2(n102), .B1(a[12]), .B2(n103), .C1(
        subAM[12]), .C2(n104), .ZN(n133) );
  INV_X1 U166 ( .A(n134), .ZN(nextA[10]) );
  AOI222_X1 U167 ( .A1(sumAM[11]), .A2(n102), .B1(a[11]), .B2(n103), .C1(
        subAM[11]), .C2(n104), .ZN(n134) );
  INV_X1 U168 ( .A(n135), .ZN(nextA[0]) );
  AOI222_X1 U169 ( .A1(sumAM[1]), .A2(n102), .B1(a[1]), .B2(n103), .C1(
        subAM[1]), .C2(n104), .ZN(n135) );
  INV_X1 U170 ( .A(q_1), .ZN(n136) );
  INV_X1 U171 ( .A(m[0]), .ZN(n64) );
  INV_X1 U172 ( .A(m[1]), .ZN(n63) );
  INV_X1 U173 ( .A(m[2]), .ZN(n62) );
  INV_X1 U174 ( .A(m[3]), .ZN(n61) );
  INV_X1 U175 ( .A(m[4]), .ZN(n60) );
  INV_X1 U176 ( .A(m[5]), .ZN(n59) );
  INV_X1 U177 ( .A(m[6]), .ZN(n58) );
  INV_X1 U178 ( .A(m[7]), .ZN(n57) );
  INV_X1 U179 ( .A(m[8]), .ZN(n56) );
  INV_X1 U180 ( .A(m[9]), .ZN(n55) );
  INV_X1 U181 ( .A(m[10]), .ZN(n54) );
  INV_X1 U182 ( .A(m[11]), .ZN(n53) );
  INV_X1 U183 ( .A(m[12]), .ZN(n52) );
  INV_X1 U184 ( .A(m[13]), .ZN(n51) );
  INV_X1 U185 ( .A(m[14]), .ZN(n50) );
  INV_X1 U186 ( .A(m[15]), .ZN(n49) );
  INV_X1 U187 ( .A(m[16]), .ZN(n48) );
  INV_X1 U188 ( .A(m[17]), .ZN(n47) );
  INV_X1 U189 ( .A(m[18]), .ZN(n46) );
  INV_X1 U190 ( .A(m[19]), .ZN(n45) );
  INV_X1 U191 ( .A(m[20]), .ZN(n44) );
  INV_X1 U192 ( .A(m[21]), .ZN(n43) );
  INV_X1 U193 ( .A(m[22]), .ZN(n42) );
  INV_X1 U194 ( .A(m[23]), .ZN(n41) );
  INV_X1 U195 ( .A(m[24]), .ZN(n40) );
  INV_X1 U196 ( .A(m[25]), .ZN(n39) );
  INV_X1 U197 ( .A(m[26]), .ZN(n38) );
  INV_X1 U198 ( .A(m[27]), .ZN(n37) );
  INV_X1 U199 ( .A(m[28]), .ZN(n36) );
  INV_X1 U200 ( .A(m[29]), .ZN(n35) );
  INV_X1 U201 ( .A(m[30]), .ZN(n34) );
  INV_X1 U202 ( .A(m[31]), .ZN(n33) );
endmodule



module regN_N32_0 ( clk, reset, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, reset;
  wire   n33, n29, n30, n31, n32, n34;

  DFF_X1 out_reg_1_ ( .D(n32), .CK(clk), .Q(out[1]) );
  DFF_X1 out_reg_0_ ( .D(n31), .CK(clk), .Q(out[0]) );
  DFF_X1 out_reg_2_ ( .D(n30), .CK(clk), .Q(out[2]) );
  DFF_X1 out_reg_5_ ( .D(n29), .CK(clk), .Q(out[5]) );
  SDFF_X1 out_reg_9_ ( .D(1'b0), .SI(n33), .SE(in[9]), .CK(clk), .Q(out[9]) );
  SDFF_X1 out_reg_8_ ( .D(1'b0), .SI(n33), .SE(in[8]), .CK(clk), .Q(out[8]) );
  SDFF_X1 out_reg_7_ ( .D(1'b0), .SI(n33), .SE(in[7]), .CK(clk), .Q(out[7]) );
  SDFF_X1 out_reg_6_ ( .D(1'b0), .SI(n33), .SE(in[6]), .CK(clk), .Q(out[6]) );
  SDFF_X1 out_reg_4_ ( .D(1'b0), .SI(n33), .SE(in[4]), .CK(clk), .Q(out[4]) );
  SDFF_X1 out_reg_3_ ( .D(1'b0), .SI(n33), .SE(in[3]), .CK(clk), .Q(out[3]) );
  SDFF_X1 out_reg_31_ ( .D(1'b0), .SI(n33), .SE(in[31]), .CK(clk), .Q(out[31])
         );
  SDFF_X1 out_reg_30_ ( .D(1'b0), .SI(n33), .SE(in[30]), .CK(clk), .Q(out[30])
         );
  SDFF_X1 out_reg_29_ ( .D(1'b0), .SI(n33), .SE(in[29]), .CK(clk), .Q(out[29])
         );
  SDFF_X1 out_reg_28_ ( .D(1'b0), .SI(n33), .SE(in[28]), .CK(clk), .Q(out[28])
         );
  SDFF_X1 out_reg_27_ ( .D(1'b0), .SI(n33), .SE(in[27]), .CK(clk), .Q(out[27])
         );
  SDFF_X1 out_reg_26_ ( .D(1'b0), .SI(n33), .SE(in[26]), .CK(clk), .Q(out[26])
         );
  SDFF_X1 out_reg_25_ ( .D(1'b0), .SI(n33), .SE(in[25]), .CK(clk), .Q(out[25])
         );
  SDFF_X1 out_reg_24_ ( .D(1'b0), .SI(n33), .SE(in[24]), .CK(clk), .Q(out[24])
         );
  SDFF_X1 out_reg_23_ ( .D(1'b0), .SI(n33), .SE(in[23]), .CK(clk), .Q(out[23])
         );
  SDFF_X1 out_reg_22_ ( .D(1'b0), .SI(n33), .SE(in[22]), .CK(clk), .Q(out[22])
         );
  SDFF_X1 out_reg_21_ ( .D(1'b0), .SI(n33), .SE(in[21]), .CK(clk), .Q(out[21])
         );
  SDFF_X1 out_reg_20_ ( .D(1'b0), .SI(n33), .SE(in[20]), .CK(clk), .Q(out[20])
         );
  SDFF_X1 out_reg_19_ ( .D(1'b0), .SI(n33), .SE(in[19]), .CK(clk), .Q(out[19])
         );
  SDFF_X1 out_reg_18_ ( .D(1'b0), .SI(n33), .SE(in[18]), .CK(clk), .Q(out[18])
         );
  SDFF_X1 out_reg_17_ ( .D(1'b0), .SI(n33), .SE(in[17]), .CK(clk), .Q(out[17])
         );
  SDFF_X1 out_reg_16_ ( .D(1'b0), .SI(n33), .SE(in[16]), .CK(clk), .Q(out[16])
         );
  SDFF_X1 out_reg_15_ ( .D(1'b0), .SI(n33), .SE(in[15]), .CK(clk), .Q(out[15])
         );
  SDFF_X1 out_reg_14_ ( .D(1'b0), .SI(n33), .SE(in[14]), .CK(clk), .Q(out[14])
         );
  SDFF_X1 out_reg_13_ ( .D(1'b0), .SI(n33), .SE(in[13]), .CK(clk), .Q(out[13])
         );
  SDFF_X1 out_reg_12_ ( .D(1'b0), .SI(n33), .SE(in[12]), .CK(clk), .Q(out[12])
         );
  SDFF_X1 out_reg_11_ ( .D(1'b0), .SI(n33), .SE(in[11]), .CK(clk), .Q(out[11])
         );
  SDFF_X1 out_reg_10_ ( .D(1'b0), .SI(n33), .SE(in[10]), .CK(clk), .Q(out[10])
         );
  BUF_X1 U31 ( .A(n33), .Z(n34) );
  INV_X1 U32 ( .A(reset), .ZN(n33) );
  AND2_X1 U33 ( .A1(in[5]), .A2(n34), .ZN(n29) );
  AND2_X1 U34 ( .A1(in[2]), .A2(n34), .ZN(n30) );
  AND2_X1 U35 ( .A1(in[0]), .A2(n34), .ZN(n31) );
  AND2_X1 U36 ( .A1(in[1]), .A2(n34), .ZN(n32) );
endmodule


module BWAdder_0 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n64, n65, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n64), .Z(result[9]) );
  XOR2_X1 U129 ( .A(n65), .B(c[8]), .Z(result[8]) );
  XOR2_X1 U131 ( .A(n67), .B(c[6]), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n68), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n68) );
  XOR2_X1 U134 ( .A(c[62]), .B(n69), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n70), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n71), .Z(result[60]) );
  XOR2_X1 U137 ( .A(n72), .B(c[5]), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n73), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n74), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n75), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n76), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n77), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n78), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n79), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n80), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n81), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n82), .Z(result[50]) );
  XOR2_X1 U148 ( .A(n83), .B(c[4]), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n84), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n85), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n86), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n87), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n88), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n89), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n90), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n91), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n92), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n93), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n94), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n95), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n96), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n97), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n98), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n99), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n100), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n101), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n102), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n103), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n104), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n105), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n106), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n107), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n108), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n109), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n110), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n111), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n112), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n113), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n114), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n115), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n116), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n117), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n118), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n119), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n120), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n121), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n122), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n123), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n124), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n125), .Z(result[11]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n127), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n65) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n67) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n72) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n69) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n70) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n71) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n73) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n83) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n74) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n75) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n76) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n77) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n78) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n79) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n80) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n81) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n82) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n84) );
  XOR2_X1 U212 ( .A(b[3]), .B(a[3]), .Z(n94) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n85) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n86) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n87) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n88) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n89) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n90) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n91) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n92) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n93) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n95) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n105) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n96) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n97) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n98) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n99) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n100) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n101) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n102) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n103) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n104) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n106) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n116) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n107) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n108) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n109) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n110) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n111) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n112) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n113) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n114) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n115) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n117) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n127) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n118) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n119) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n120) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n121) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n122) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n123) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n124) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n125) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n126) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n64) );
  CLKBUF_X1 U2 ( .A(n65), .Z(n1) );
  CLKBUF_X1 U3 ( .A(b[5]), .Z(n2) );
  XNOR2_X1 U4 ( .A(n3), .B(c[7]), .ZN(result[7]) );
  XNOR2_X1 U5 ( .A(a[7]), .B(b[7]), .ZN(n3) );
  CLKBUF_X1 U6 ( .A(b[8]), .Z(n4) );
  CLKBUF_X1 U7 ( .A(a[8]), .Z(n5) );
  NAND2_X1 U8 ( .A1(c[10]), .A2(n7), .ZN(n8) );
  NAND2_X1 U9 ( .A1(n6), .A2(n126), .ZN(n9) );
  NAND2_X1 U10 ( .A1(n8), .A2(n9), .ZN(result[10]) );
  INV_X1 U11 ( .A(c[10]), .ZN(n6) );
  INV_X1 U12 ( .A(n126), .ZN(n7) );
  XOR2_X1 U13 ( .A(a[7]), .B(b[7]), .Z(n10) );
  INV_X1 U14 ( .A(n158), .ZN(carry[3]) );
  AOI22_X1 U15 ( .A1(b[2]), .A2(a[2]), .B1(n105), .B2(c[2]), .ZN(n158) );
  INV_X1 U16 ( .A(n182), .ZN(carry[18]) );
  AOI22_X1 U17 ( .A1(b[17]), .A2(a[17]), .B1(n119), .B2(c[17]), .ZN(n182) );
  INV_X1 U18 ( .A(n181), .ZN(carry[19]) );
  AOI22_X1 U19 ( .A1(b[18]), .A2(a[18]), .B1(n118), .B2(c[18]), .ZN(n181) );
  INV_X1 U20 ( .A(n189), .ZN(carry[11]) );
  AOI22_X1 U21 ( .A1(b[10]), .A2(a[10]), .B1(n126), .B2(c[10]), .ZN(n189) );
  INV_X1 U22 ( .A(n186), .ZN(carry[14]) );
  AOI22_X1 U23 ( .A1(b[13]), .A2(a[13]), .B1(n123), .B2(c[13]), .ZN(n186) );
  INV_X1 U24 ( .A(n179), .ZN(carry[20]) );
  AOI22_X1 U25 ( .A1(b[19]), .A2(a[19]), .B1(n117), .B2(c[19]), .ZN(n179) );
  INV_X1 U26 ( .A(n178), .ZN(carry[21]) );
  AOI22_X1 U27 ( .A1(b[20]), .A2(a[20]), .B1(n115), .B2(c[20]), .ZN(n178) );
  INV_X1 U28 ( .A(n177), .ZN(carry[22]) );
  AOI22_X1 U29 ( .A1(b[21]), .A2(a[21]), .B1(n114), .B2(c[21]), .ZN(n177) );
  INV_X1 U30 ( .A(n176), .ZN(carry[23]) );
  AOI22_X1 U31 ( .A1(b[22]), .A2(a[22]), .B1(n113), .B2(c[22]), .ZN(n176) );
  INV_X1 U32 ( .A(n147), .ZN(carry[4]) );
  INV_X1 U33 ( .A(n183), .ZN(carry[17]) );
  AOI22_X1 U34 ( .A1(b[16]), .A2(a[16]), .B1(n120), .B2(c[16]), .ZN(n183) );
  INV_X1 U35 ( .A(n188), .ZN(carry[12]) );
  AOI22_X1 U36 ( .A1(b[11]), .A2(a[11]), .B1(n125), .B2(c[11]), .ZN(n188) );
  INV_X1 U37 ( .A(n187), .ZN(carry[13]) );
  AOI22_X1 U38 ( .A1(b[12]), .A2(a[12]), .B1(n124), .B2(c[12]), .ZN(n187) );
  INV_X1 U39 ( .A(n185), .ZN(carry[15]) );
  AOI22_X1 U40 ( .A1(b[14]), .A2(a[14]), .B1(n122), .B2(c[14]), .ZN(n185) );
  INV_X1 U41 ( .A(n184), .ZN(carry[16]) );
  AOI22_X1 U42 ( .A1(b[15]), .A2(a[15]), .B1(n121), .B2(c[15]), .ZN(n184) );
  INV_X1 U43 ( .A(n175), .ZN(carry[24]) );
  AOI22_X1 U44 ( .A1(b[23]), .A2(a[23]), .B1(n112), .B2(c[23]), .ZN(n175) );
  INV_X1 U45 ( .A(n174), .ZN(carry[25]) );
  AOI22_X1 U46 ( .A1(b[24]), .A2(a[24]), .B1(n111), .B2(c[24]), .ZN(n174) );
  INV_X1 U47 ( .A(n173), .ZN(carry[26]) );
  AOI22_X1 U48 ( .A1(b[25]), .A2(a[25]), .B1(n110), .B2(c[25]), .ZN(n173) );
  INV_X1 U49 ( .A(n172), .ZN(carry[27]) );
  AOI22_X1 U50 ( .A1(b[26]), .A2(a[26]), .B1(n109), .B2(c[26]), .ZN(n172) );
  INV_X1 U51 ( .A(n171), .ZN(carry[28]) );
  AOI22_X1 U52 ( .A1(b[27]), .A2(a[27]), .B1(n108), .B2(c[27]), .ZN(n171) );
  INV_X1 U53 ( .A(n170), .ZN(carry[29]) );
  AOI22_X1 U54 ( .A1(b[28]), .A2(a[28]), .B1(n107), .B2(c[28]), .ZN(n170) );
  INV_X1 U55 ( .A(n168), .ZN(carry[30]) );
  AOI22_X1 U56 ( .A1(b[29]), .A2(a[29]), .B1(n106), .B2(c[29]), .ZN(n168) );
  INV_X1 U57 ( .A(n190), .ZN(carry[10]) );
  AOI22_X1 U58 ( .A1(b[9]), .A2(a[9]), .B1(n64), .B2(c[9]), .ZN(n190) );
  INV_X1 U59 ( .A(n136), .ZN(carry[5]) );
  INV_X1 U60 ( .A(n130), .ZN(carry[7]) );
  INV_X1 U61 ( .A(n131), .ZN(carry[6]) );
  INV_X1 U62 ( .A(n129), .ZN(carry[8]) );
  INV_X1 U63 ( .A(n128), .ZN(carry[9]) );
  INV_X1 U64 ( .A(n161), .ZN(carry[37]) );
  AOI22_X1 U65 ( .A1(b[36]), .A2(a[36]), .B1(n98), .B2(c[36]), .ZN(n161) );
  INV_X1 U66 ( .A(n160), .ZN(carry[38]) );
  AOI22_X1 U67 ( .A1(b[37]), .A2(a[37]), .B1(n97), .B2(c[37]), .ZN(n160) );
  INV_X1 U68 ( .A(n159), .ZN(carry[39]) );
  AOI22_X1 U69 ( .A1(b[38]), .A2(a[38]), .B1(n96), .B2(c[38]), .ZN(n159) );
  INV_X1 U70 ( .A(n157), .ZN(carry[40]) );
  AOI22_X1 U71 ( .A1(b[39]), .A2(a[39]), .B1(n95), .B2(c[39]), .ZN(n157) );
  INV_X1 U72 ( .A(n156), .ZN(carry[41]) );
  AOI22_X1 U73 ( .A1(b[40]), .A2(a[40]), .B1(n93), .B2(c[40]), .ZN(n156) );
  INV_X1 U74 ( .A(n155), .ZN(carry[42]) );
  AOI22_X1 U75 ( .A1(b[41]), .A2(a[41]), .B1(n92), .B2(c[41]), .ZN(n155) );
  INV_X1 U76 ( .A(n165), .ZN(carry[33]) );
  AOI22_X1 U77 ( .A1(b[32]), .A2(a[32]), .B1(n102), .B2(c[32]), .ZN(n165) );
  INV_X1 U78 ( .A(n164), .ZN(carry[34]) );
  AOI22_X1 U79 ( .A1(b[33]), .A2(a[33]), .B1(n101), .B2(c[33]), .ZN(n164) );
  INV_X1 U80 ( .A(n163), .ZN(carry[35]) );
  AOI22_X1 U81 ( .A1(b[34]), .A2(a[34]), .B1(n100), .B2(c[34]), .ZN(n163) );
  INV_X1 U82 ( .A(n162), .ZN(carry[36]) );
  AOI22_X1 U83 ( .A1(b[35]), .A2(a[35]), .B1(n99), .B2(c[35]), .ZN(n162) );
  INV_X1 U84 ( .A(n167), .ZN(carry[31]) );
  AOI22_X1 U85 ( .A1(b[30]), .A2(a[30]), .B1(n104), .B2(c[30]), .ZN(n167) );
  INV_X1 U86 ( .A(n166), .ZN(carry[32]) );
  AOI22_X1 U87 ( .A1(b[31]), .A2(a[31]), .B1(n103), .B2(c[31]), .ZN(n166) );
  INV_X1 U88 ( .A(n154), .ZN(carry[43]) );
  AOI22_X1 U89 ( .A1(b[42]), .A2(a[42]), .B1(n91), .B2(c[42]), .ZN(n154) );
  INV_X1 U90 ( .A(n153), .ZN(carry[44]) );
  AOI22_X1 U91 ( .A1(b[43]), .A2(a[43]), .B1(n90), .B2(c[43]), .ZN(n153) );
  INV_X1 U92 ( .A(n152), .ZN(carry[45]) );
  AOI22_X1 U93 ( .A1(b[44]), .A2(a[44]), .B1(n89), .B2(c[44]), .ZN(n152) );
  INV_X1 U94 ( .A(n151), .ZN(carry[46]) );
  AOI22_X1 U95 ( .A1(b[45]), .A2(a[45]), .B1(n88), .B2(c[45]), .ZN(n151) );
  INV_X1 U96 ( .A(n150), .ZN(carry[47]) );
  AOI22_X1 U97 ( .A1(b[46]), .A2(a[46]), .B1(n87), .B2(c[46]), .ZN(n150) );
  INV_X1 U98 ( .A(n149), .ZN(carry[48]) );
  AOI22_X1 U99 ( .A1(b[47]), .A2(a[47]), .B1(n86), .B2(c[47]), .ZN(n149) );
  INV_X1 U100 ( .A(n148), .ZN(carry[49]) );
  AOI22_X1 U101 ( .A1(b[48]), .A2(a[48]), .B1(n85), .B2(c[48]), .ZN(n148) );
  INV_X1 U102 ( .A(n146), .ZN(carry[50]) );
  AOI22_X1 U103 ( .A1(b[49]), .A2(a[49]), .B1(n84), .B2(c[49]), .ZN(n146) );
  INV_X1 U104 ( .A(n145), .ZN(carry[51]) );
  AOI22_X1 U105 ( .A1(b[50]), .A2(a[50]), .B1(n82), .B2(c[50]), .ZN(n145) );
  INV_X1 U106 ( .A(n144), .ZN(carry[52]) );
  AOI22_X1 U107 ( .A1(b[51]), .A2(a[51]), .B1(n81), .B2(c[51]), .ZN(n144) );
  INV_X1 U108 ( .A(n143), .ZN(carry[53]) );
  AOI22_X1 U109 ( .A1(b[52]), .A2(a[52]), .B1(n80), .B2(c[52]), .ZN(n143) );
  INV_X1 U110 ( .A(n142), .ZN(carry[54]) );
  AOI22_X1 U111 ( .A1(b[53]), .A2(a[53]), .B1(n79), .B2(c[53]), .ZN(n142) );
  INV_X1 U112 ( .A(n141), .ZN(carry[55]) );
  AOI22_X1 U113 ( .A1(b[54]), .A2(a[54]), .B1(n78), .B2(c[54]), .ZN(n141) );
  INV_X1 U114 ( .A(n140), .ZN(carry[56]) );
  AOI22_X1 U115 ( .A1(b[55]), .A2(a[55]), .B1(n77), .B2(c[55]), .ZN(n140) );
  INV_X1 U116 ( .A(n139), .ZN(carry[57]) );
  AOI22_X1 U117 ( .A1(b[56]), .A2(a[56]), .B1(n76), .B2(c[56]), .ZN(n139) );
  INV_X1 U118 ( .A(n138), .ZN(carry[58]) );
  AOI22_X1 U119 ( .A1(b[57]), .A2(a[57]), .B1(n75), .B2(c[57]), .ZN(n138) );
  INV_X1 U120 ( .A(n137), .ZN(carry[59]) );
  AOI22_X1 U121 ( .A1(b[58]), .A2(a[58]), .B1(n74), .B2(c[58]), .ZN(n137) );
  INV_X1 U122 ( .A(n135), .ZN(carry[60]) );
  AOI22_X1 U123 ( .A1(b[59]), .A2(a[59]), .B1(n73), .B2(c[59]), .ZN(n135) );
  INV_X1 U124 ( .A(n134), .ZN(carry[61]) );
  AOI22_X1 U125 ( .A1(b[60]), .A2(a[60]), .B1(n71), .B2(c[60]), .ZN(n134) );
  INV_X1 U126 ( .A(n133), .ZN(carry[62]) );
  AOI22_X1 U127 ( .A1(b[61]), .A2(a[61]), .B1(n70), .B2(c[61]), .ZN(n133) );
  INV_X1 U130 ( .A(n132), .ZN(carry[63]) );
  AOI22_X1 U191 ( .A1(b[62]), .A2(a[62]), .B1(n69), .B2(c[62]), .ZN(n132) );
  INV_X1 U194 ( .A(n169), .ZN(carry[2]) );
  AOI22_X1 U256 ( .A1(b[1]), .A2(a[1]), .B1(n116), .B2(c[1]), .ZN(n169) );
  INV_X1 U257 ( .A(n180), .ZN(carry[1]) );
  AOI22_X1 U258 ( .A1(b[0]), .A2(a[0]), .B1(n127), .B2(c[0]), .ZN(n180) );
  AOI22_X1 U259 ( .A1(b[3]), .A2(a[3]), .B1(n94), .B2(c[3]), .ZN(n147) );
  CLKBUF_X1 U260 ( .A(a[5]), .Z(n11) );
  AOI22_X1 U261 ( .A1(b[4]), .A2(a[4]), .B1(n83), .B2(c[4]), .ZN(n136) );
  AOI22_X1 U262 ( .A1(b[6]), .A2(a[6]), .B1(n67), .B2(c[6]), .ZN(n130) );
  AOI22_X1 U263 ( .A1(n4), .A2(n5), .B1(n1), .B2(c[8]), .ZN(n128) );
  AOI22_X1 U264 ( .A1(n2), .A2(n11), .B1(n72), .B2(c[5]), .ZN(n131) );
  AOI22_X1 U265 ( .A1(b[7]), .A2(a[7]), .B1(n10), .B2(c[7]), .ZN(n129) );
endmodule


module FullAdder_0 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(cin), .B(n2), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(cout) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(n2), .B2(cin), .ZN(n3) );
endmodule


module FullAdder_1 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5, n6;

  XOR2_X1 U4 ( .A(a), .B(b), .Z(n6) );
  INV_X1 U1 ( .A(n6), .ZN(n4) );
  CLKBUF_X1 U2 ( .A(cin), .Z(n1) );
  XNOR2_X1 U3 ( .A(cin), .B(n4), .ZN(sum) );
  INV_X1 U5 ( .A(n5), .ZN(cout) );
  AOI22_X1 U6 ( .A1(b), .A2(a), .B1(n6), .B2(n1), .ZN(n5) );
endmodule


module FullAdder_2 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_3 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(cin), .B(n3), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(cout) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n3), .ZN(n1) );
endmodule


module FullAdder_4 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_5 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(cin), .B(n3), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(cout) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n3), .ZN(n1) );
endmodule


module FullAdder_6 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(cin), .B(n3), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(cout) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n3), .ZN(n1) );
endmodule


module FullAdder_7 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_8 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_9 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_10 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_11 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_12 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_13 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_14 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_15 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_16 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_17 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_18 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_19 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_20 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_21 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_22 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_23 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_24 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  XOR2_X1 U2 ( .A(n1), .B(n5), .Z(sum) );
  INV_X1 U3 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_25 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_26 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_27 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_28 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_29 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_30 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(cin), .B(n3), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n3) );
  AOI22_X1 U1 ( .A1(b), .A2(a), .B1(cin), .B2(n3), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(cout) );
endmodule


module FullAdder_31 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_32 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_33 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_34 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_35 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_36 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(cin), .B(n3), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(cout) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n3), .ZN(n1) );
endmodule


module FullAdder_37 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_38 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_39 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_40 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(cin), .B(n3), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n3) );
  AOI22_X1 U1 ( .A1(b), .A2(a), .B1(cin), .B2(n3), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(cout) );
endmodule


module FullAdder_41 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_42 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_43 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_44 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_45 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_46 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_47 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_48 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_49 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_50 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_51 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_52 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(n1), .B(n5), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(cin), .Z(n1) );
  INV_X1 U2 ( .A(n4), .ZN(cout) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
endmodule


module FullAdder_53 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5;

  XOR2_X1 U3 ( .A(cin), .B(n1), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n5) );
  CLKBUF_X1 U1 ( .A(n5), .Z(n1) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(cin), .B2(n5), .ZN(n4) );
  INV_X1 U5 ( .A(n4), .ZN(cout) );
endmodule


module FullAdder_54 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5, n6;

  XOR2_X1 U3 ( .A(n4), .B(n1), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n6) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n1) );
  CLKBUF_X1 U2 ( .A(cin), .Z(n4) );
  AOI22_X1 U5 ( .A1(b), .A2(a), .B1(cin), .B2(n6), .ZN(n5) );
  INV_X1 U6 ( .A(n5), .ZN(cout) );
endmodule


module FullAdder_55 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5, n6;

  XOR2_X1 U3 ( .A(cin), .B(n4), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n6) );
  CLKBUF_X1 U1 ( .A(a), .Z(n1) );
  CLKBUF_X1 U2 ( .A(n6), .Z(n4) );
  AOI22_X1 U5 ( .A1(b), .A2(n1), .B1(cin), .B2(n6), .ZN(n5) );
  INV_X1 U6 ( .A(n5), .ZN(cout) );
endmodule


module FullAdder_56 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n4, n5, n6;

  XOR2_X1 U3 ( .A(cin), .B(n4), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n6) );
  CLKBUF_X1 U1 ( .A(a), .Z(n1) );
  CLKBUF_X1 U2 ( .A(n6), .Z(n4) );
  AOI22_X1 U5 ( .A1(b), .A2(n1), .B1(n6), .B2(cin), .ZN(n5) );
  INV_X1 U6 ( .A(n5), .ZN(cout) );
endmodule


module FullAdder_57 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(cin), .B(n3), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n3) );
  AOI22_X1 U1 ( .A1(b), .A2(a), .B1(n3), .B2(cin), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(cout) );
endmodule


module FullAdder_58 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(cin), .B(n3), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n3) );
  AOI22_X1 U1 ( .A1(b), .A2(a), .B1(n3), .B2(cin), .ZN(n1) );
  INV_X1 U2 ( .A(n1), .ZN(cout) );
endmodule


module FullAdder_59 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(cin), .B(n3), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(cout) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(n3), .B2(cin), .ZN(n1) );
endmodule


module FullAdder_60 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(cin), .B(n3), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(cout) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(n3), .B2(cin), .ZN(n1) );
endmodule


module FullAdder_61 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(cin), .B(n3), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(cout) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(n3), .B2(cin), .ZN(n1) );
endmodule


module FullAdder_62 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(cin), .B(n3), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(cout) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(n3), .B2(cin), .ZN(n1) );
endmodule


module FullAdder_63 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n3;

  XOR2_X1 U3 ( .A(cin), .B(n3), .Z(sum) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n3) );
  INV_X1 U1 ( .A(n1), .ZN(cout) );
  AOI22_X1 U2 ( .A1(b), .A2(a), .B1(n3), .B2(cin), .ZN(n1) );
endmodule


module CRAdder_64 ( a, b, cin, sum, cout, overflow );
  input [63:0] a;
  input [63:0] b;
  output [63:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2, n3;
  wire   [62:0] passCout;

  FullAdder_0 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_63 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_62 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_61 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_60 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_59 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_58 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_57 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_56 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_55 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_54 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_53 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_52 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_51 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_50 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_49 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_48 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_47 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_46 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_45 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_44 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_43 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_42 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_41 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_40 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_39 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_38 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_37 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_36 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_35 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_34 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_33 bit_gen_31__bit ( .a(a[31]), .b(b[31]), .cin(passCout[30]), 
        .sum(sum[31]), .cout(passCout[31]) );
  FullAdder_32 bit_gen_32__bit ( .a(a[32]), .b(b[32]), .cin(passCout[31]), 
        .sum(sum[32]), .cout(passCout[32]) );
  FullAdder_31 bit_gen_33__bit ( .a(a[33]), .b(b[33]), .cin(passCout[32]), 
        .sum(sum[33]), .cout(passCout[33]) );
  FullAdder_30 bit_gen_34__bit ( .a(a[34]), .b(b[34]), .cin(passCout[33]), 
        .sum(sum[34]), .cout(passCout[34]) );
  FullAdder_29 bit_gen_35__bit ( .a(a[35]), .b(b[35]), .cin(passCout[34]), 
        .sum(sum[35]), .cout(passCout[35]) );
  FullAdder_28 bit_gen_36__bit ( .a(a[36]), .b(b[36]), .cin(passCout[35]), 
        .sum(sum[36]), .cout(passCout[36]) );
  FullAdder_27 bit_gen_37__bit ( .a(a[37]), .b(b[37]), .cin(passCout[36]), 
        .sum(sum[37]), .cout(passCout[37]) );
  FullAdder_26 bit_gen_38__bit ( .a(a[38]), .b(b[38]), .cin(passCout[37]), 
        .sum(sum[38]), .cout(passCout[38]) );
  FullAdder_25 bit_gen_39__bit ( .a(a[39]), .b(b[39]), .cin(passCout[38]), 
        .sum(sum[39]), .cout(passCout[39]) );
  FullAdder_24 bit_gen_40__bit ( .a(a[40]), .b(b[40]), .cin(passCout[39]), 
        .sum(sum[40]), .cout(passCout[40]) );
  FullAdder_23 bit_gen_41__bit ( .a(a[41]), .b(b[41]), .cin(passCout[40]), 
        .sum(sum[41]), .cout(passCout[41]) );
  FullAdder_22 bit_gen_42__bit ( .a(a[42]), .b(b[42]), .cin(passCout[41]), 
        .sum(sum[42]), .cout(passCout[42]) );
  FullAdder_21 bit_gen_43__bit ( .a(a[43]), .b(b[43]), .cin(passCout[42]), 
        .sum(sum[43]), .cout(passCout[43]) );
  FullAdder_20 bit_gen_44__bit ( .a(a[44]), .b(b[44]), .cin(passCout[43]), 
        .sum(sum[44]), .cout(passCout[44]) );
  FullAdder_19 bit_gen_45__bit ( .a(a[45]), .b(b[45]), .cin(passCout[44]), 
        .sum(sum[45]), .cout(passCout[45]) );
  FullAdder_18 bit_gen_46__bit ( .a(a[46]), .b(b[46]), .cin(passCout[45]), 
        .sum(sum[46]), .cout(passCout[46]) );
  FullAdder_17 bit_gen_47__bit ( .a(a[47]), .b(b[47]), .cin(passCout[46]), 
        .sum(sum[47]), .cout(passCout[47]) );
  FullAdder_16 bit_gen_48__bit ( .a(a[48]), .b(b[48]), .cin(passCout[47]), 
        .sum(sum[48]), .cout(passCout[48]) );
  FullAdder_15 bit_gen_49__bit ( .a(a[49]), .b(b[49]), .cin(passCout[48]), 
        .sum(sum[49]), .cout(passCout[49]) );
  FullAdder_14 bit_gen_50__bit ( .a(a[50]), .b(b[50]), .cin(passCout[49]), 
        .sum(sum[50]), .cout(passCout[50]) );
  FullAdder_13 bit_gen_51__bit ( .a(a[51]), .b(b[51]), .cin(passCout[50]), 
        .sum(sum[51]), .cout(passCout[51]) );
  FullAdder_12 bit_gen_52__bit ( .a(a[52]), .b(b[52]), .cin(passCout[51]), 
        .sum(sum[52]), .cout(passCout[52]) );
  FullAdder_11 bit_gen_53__bit ( .a(a[53]), .b(b[53]), .cin(passCout[52]), 
        .sum(sum[53]), .cout(passCout[53]) );
  FullAdder_10 bit_gen_54__bit ( .a(a[54]), .b(b[54]), .cin(passCout[53]), 
        .sum(sum[54]), .cout(passCout[54]) );
  FullAdder_9 bit_gen_55__bit ( .a(a[55]), .b(b[55]), .cin(passCout[54]), 
        .sum(sum[55]), .cout(passCout[55]) );
  FullAdder_8 bit_gen_56__bit ( .a(a[56]), .b(b[56]), .cin(passCout[55]), 
        .sum(sum[56]), .cout(passCout[56]) );
  FullAdder_7 bit_gen_57__bit ( .a(a[57]), .b(b[57]), .cin(passCout[56]), 
        .sum(sum[57]), .cout(passCout[57]) );
  FullAdder_6 bit_gen_58__bit ( .a(a[58]), .b(b[58]), .cin(passCout[57]), 
        .sum(sum[58]), .cout(passCout[58]) );
  FullAdder_5 bit_gen_59__bit ( .a(a[59]), .b(b[59]), .cin(passCout[58]), 
        .sum(sum[59]), .cout(passCout[59]) );
  FullAdder_4 bit_gen_60__bit ( .a(a[60]), .b(b[60]), .cin(passCout[59]), 
        .sum(sum[60]), .cout(passCout[60]) );
  FullAdder_3 bit_gen_61__bit ( .a(a[61]), .b(b[61]), .cin(passCout[60]), 
        .sum(sum[61]), .cout(passCout[61]) );
  FullAdder_2 bit_gen_62__bit ( .a(a[62]), .b(b[62]), .cin(passCout[61]), 
        .sum(sum[62]), .cout(passCout[62]) );
  FullAdder_1 bit63 ( .a(a[63]), .b(b[63]), .cin(passCout[62]), .sum(sum[63]), 
        .cout(cout) );
  XOR2_X1 U3 ( .A(b[63]), .B(a[63]), .Z(n2) );
  CLKBUF_X1 U1 ( .A(sum[63]), .Z(n3) );
  XNOR2_X1 U2 ( .A(a[63]), .B(n3), .ZN(n1) );
  NOR2_X1 U4 ( .A1(n1), .A2(n2), .ZN(overflow) );
endmodule


module BWAdder_1 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(n213), .B(c[9]), .Z(result[9]) );
  XOR2_X1 U129 ( .A(n212), .B(c[8]), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n211), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n209), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n209) );
  XOR2_X1 U134 ( .A(c[62]), .B(n208), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n207), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n206), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n205), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n204), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n203), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n202), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n201), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n200), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n199), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n198), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n197), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n196), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n195), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n194), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n193), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n192), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n191), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n190), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n189), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n188), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n187), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n186), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n185), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n184), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n183), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n182), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n181), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n180), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n179), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n178), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n177), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n176), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n175), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n174), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n173), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n172), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n171), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n170), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n169), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n168), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n167), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n166), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n165), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n164), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n163), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n162), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n161), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n160), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n159), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n158), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n157), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n156), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n155), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n154), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n153), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n152), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n151), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n150), .Z(result[0]) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n205) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n208) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n207) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n206) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n204) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n194) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n203) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n202) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n201) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n200) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n199) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n198) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n197) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n196) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n195) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n193) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n183) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n192) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n191) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n190) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n189) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n188) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n187) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n186) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n185) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n184) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n182) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n172) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n181) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n180) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n179) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n178) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n177) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n176) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n175) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n174) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n173) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n171) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n161) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n170) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n169) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n168) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n167) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n166) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n165) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n164) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n163) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n162) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n160) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n150) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n159) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n158) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n157) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n156) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n155) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n154) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n153) );
  INV_X1 U2 ( .A(b[11]), .ZN(n3) );
  INV_X1 U3 ( .A(b[10]), .ZN(n5) );
  INV_X1 U4 ( .A(b[9]), .ZN(n10) );
  INV_X1 U5 ( .A(b[7]), .ZN(n9) );
  INV_X1 U6 ( .A(b[6]), .ZN(n8) );
  CLKBUF_X1 U7 ( .A(a[6]), .Z(n1) );
  CLKBUF_X1 U8 ( .A(a[8]), .Z(n2) );
  XNOR2_X1 U9 ( .A(a[11]), .B(n3), .ZN(n152) );
  CLKBUF_X1 U10 ( .A(n210), .Z(n4) );
  XNOR2_X1 U11 ( .A(a[10]), .B(n5), .ZN(n151) );
  CLKBUF_X1 U12 ( .A(n212), .Z(n6) );
  CLKBUF_X1 U13 ( .A(a[7]), .Z(n7) );
  XNOR2_X1 U14 ( .A(a[6]), .B(n8), .ZN(n210) );
  XNOR2_X1 U15 ( .A(a[7]), .B(n9), .ZN(n211) );
  XNOR2_X1 U16 ( .A(a[9]), .B(n10), .ZN(n213) );
  INV_X1 U17 ( .A(b[8]), .ZN(n11) );
  XNOR2_X1 U18 ( .A(a[8]), .B(n11), .ZN(n212) );
  INV_X1 U19 ( .A(n149), .ZN(carry[9]) );
  INV_X1 U20 ( .A(n12), .ZN(carry[10]) );
  INV_X1 U21 ( .A(n13), .ZN(carry[11]) );
  INV_X1 U22 ( .A(n25), .ZN(carry[22]) );
  AOI22_X1 U23 ( .A1(b[21]), .A2(a[21]), .B1(n163), .B2(c[21]), .ZN(n25) );
  INV_X1 U24 ( .A(n24), .ZN(carry[21]) );
  AOI22_X1 U25 ( .A1(b[20]), .A2(a[20]), .B1(n162), .B2(c[20]), .ZN(n24) );
  INV_X1 U26 ( .A(n23), .ZN(carry[20]) );
  AOI22_X1 U27 ( .A1(b[19]), .A2(a[19]), .B1(n160), .B2(c[19]), .ZN(n23) );
  INV_X1 U28 ( .A(n14), .ZN(carry[12]) );
  AOI22_X1 U29 ( .A1(b[11]), .A2(a[11]), .B1(n152), .B2(c[11]), .ZN(n14) );
  INV_X1 U30 ( .A(n15), .ZN(carry[13]) );
  AOI22_X1 U31 ( .A1(b[12]), .A2(a[12]), .B1(n153), .B2(c[12]), .ZN(n15) );
  INV_X1 U32 ( .A(n16), .ZN(carry[14]) );
  AOI22_X1 U33 ( .A1(b[13]), .A2(a[13]), .B1(n154), .B2(c[13]), .ZN(n16) );
  INV_X1 U34 ( .A(n20), .ZN(carry[18]) );
  AOI22_X1 U35 ( .A1(b[17]), .A2(a[17]), .B1(n158), .B2(c[17]), .ZN(n20) );
  INV_X1 U36 ( .A(n17), .ZN(carry[15]) );
  AOI22_X1 U37 ( .A1(b[14]), .A2(a[14]), .B1(n155), .B2(c[14]), .ZN(n17) );
  INV_X1 U38 ( .A(n18), .ZN(carry[16]) );
  AOI22_X1 U39 ( .A1(b[15]), .A2(a[15]), .B1(n156), .B2(c[15]), .ZN(n18) );
  INV_X1 U40 ( .A(n21), .ZN(carry[19]) );
  AOI22_X1 U41 ( .A1(b[18]), .A2(a[18]), .B1(n159), .B2(c[18]), .ZN(n21) );
  INV_X1 U42 ( .A(n19), .ZN(carry[17]) );
  AOI22_X1 U43 ( .A1(b[16]), .A2(a[16]), .B1(n157), .B2(c[16]), .ZN(n19) );
  INV_X1 U44 ( .A(n26), .ZN(carry[23]) );
  AOI22_X1 U45 ( .A1(b[22]), .A2(a[22]), .B1(n164), .B2(c[22]), .ZN(n26) );
  INV_X1 U46 ( .A(n27), .ZN(carry[24]) );
  AOI22_X1 U47 ( .A1(b[23]), .A2(a[23]), .B1(n165), .B2(c[23]), .ZN(n27) );
  INV_X1 U48 ( .A(n28), .ZN(carry[25]) );
  AOI22_X1 U49 ( .A1(b[24]), .A2(a[24]), .B1(n166), .B2(c[24]), .ZN(n28) );
  INV_X1 U50 ( .A(n29), .ZN(carry[26]) );
  AOI22_X1 U51 ( .A1(b[25]), .A2(a[25]), .B1(n167), .B2(c[25]), .ZN(n29) );
  INV_X1 U52 ( .A(n30), .ZN(carry[27]) );
  AOI22_X1 U53 ( .A1(b[26]), .A2(a[26]), .B1(n168), .B2(c[26]), .ZN(n30) );
  INV_X1 U54 ( .A(n31), .ZN(carry[28]) );
  AOI22_X1 U55 ( .A1(b[27]), .A2(a[27]), .B1(n169), .B2(c[27]), .ZN(n31) );
  INV_X1 U56 ( .A(n32), .ZN(carry[29]) );
  AOI22_X1 U57 ( .A1(b[28]), .A2(a[28]), .B1(n170), .B2(c[28]), .ZN(n32) );
  INV_X1 U58 ( .A(n34), .ZN(carry[30]) );
  AOI22_X1 U59 ( .A1(b[29]), .A2(a[29]), .B1(n171), .B2(c[29]), .ZN(n34) );
  INV_X1 U60 ( .A(n35), .ZN(carry[31]) );
  AOI22_X1 U61 ( .A1(b[30]), .A2(a[30]), .B1(n173), .B2(c[30]), .ZN(n35) );
  INV_X1 U62 ( .A(n36), .ZN(carry[32]) );
  AOI22_X1 U63 ( .A1(b[31]), .A2(a[31]), .B1(n174), .B2(c[31]), .ZN(n36) );
  INV_X1 U64 ( .A(n37), .ZN(carry[33]) );
  AOI22_X1 U65 ( .A1(b[32]), .A2(a[32]), .B1(n175), .B2(c[32]), .ZN(n37) );
  INV_X1 U66 ( .A(n38), .ZN(carry[34]) );
  AOI22_X1 U67 ( .A1(b[33]), .A2(a[33]), .B1(n176), .B2(c[33]), .ZN(n38) );
  INV_X1 U68 ( .A(n39), .ZN(carry[35]) );
  AOI22_X1 U69 ( .A1(b[34]), .A2(a[34]), .B1(n177), .B2(c[34]), .ZN(n39) );
  INV_X1 U70 ( .A(n40), .ZN(carry[36]) );
  AOI22_X1 U71 ( .A1(b[35]), .A2(a[35]), .B1(n178), .B2(c[35]), .ZN(n40) );
  INV_X1 U72 ( .A(n41), .ZN(carry[37]) );
  AOI22_X1 U73 ( .A1(b[36]), .A2(a[36]), .B1(n179), .B2(c[36]), .ZN(n41) );
  INV_X1 U74 ( .A(n42), .ZN(carry[38]) );
  AOI22_X1 U75 ( .A1(b[37]), .A2(a[37]), .B1(n180), .B2(c[37]), .ZN(n42) );
  INV_X1 U76 ( .A(n43), .ZN(carry[39]) );
  AOI22_X1 U77 ( .A1(b[38]), .A2(a[38]), .B1(n181), .B2(c[38]), .ZN(n43) );
  INV_X1 U78 ( .A(n45), .ZN(carry[40]) );
  AOI22_X1 U79 ( .A1(b[39]), .A2(a[39]), .B1(n182), .B2(c[39]), .ZN(n45) );
  INV_X1 U80 ( .A(n46), .ZN(carry[41]) );
  AOI22_X1 U81 ( .A1(b[40]), .A2(a[40]), .B1(n184), .B2(c[40]), .ZN(n46) );
  INV_X1 U82 ( .A(n47), .ZN(carry[42]) );
  AOI22_X1 U83 ( .A1(b[41]), .A2(a[41]), .B1(n185), .B2(c[41]), .ZN(n47) );
  INV_X1 U84 ( .A(n48), .ZN(carry[43]) );
  AOI22_X1 U85 ( .A1(b[42]), .A2(a[42]), .B1(n186), .B2(c[42]), .ZN(n48) );
  INV_X1 U86 ( .A(n49), .ZN(carry[44]) );
  AOI22_X1 U87 ( .A1(b[43]), .A2(a[43]), .B1(n187), .B2(c[43]), .ZN(n49) );
  INV_X1 U88 ( .A(n57), .ZN(carry[51]) );
  AOI22_X1 U89 ( .A1(b[50]), .A2(a[50]), .B1(n195), .B2(c[50]), .ZN(n57) );
  INV_X1 U90 ( .A(n50), .ZN(carry[45]) );
  AOI22_X1 U91 ( .A1(b[44]), .A2(a[44]), .B1(n188), .B2(c[44]), .ZN(n50) );
  INV_X1 U92 ( .A(n51), .ZN(carry[46]) );
  AOI22_X1 U93 ( .A1(b[45]), .A2(a[45]), .B1(n189), .B2(c[45]), .ZN(n51) );
  INV_X1 U94 ( .A(n52), .ZN(carry[47]) );
  AOI22_X1 U95 ( .A1(b[46]), .A2(a[46]), .B1(n190), .B2(c[46]), .ZN(n52) );
  INV_X1 U96 ( .A(n53), .ZN(carry[48]) );
  AOI22_X1 U97 ( .A1(b[47]), .A2(a[47]), .B1(n191), .B2(c[47]), .ZN(n53) );
  INV_X1 U98 ( .A(n54), .ZN(carry[49]) );
  AOI22_X1 U99 ( .A1(b[48]), .A2(a[48]), .B1(n192), .B2(c[48]), .ZN(n54) );
  INV_X1 U100 ( .A(n56), .ZN(carry[50]) );
  AOI22_X1 U101 ( .A1(b[49]), .A2(a[49]), .B1(n193), .B2(c[49]), .ZN(n56) );
  INV_X1 U102 ( .A(n58), .ZN(carry[52]) );
  AOI22_X1 U103 ( .A1(b[51]), .A2(a[51]), .B1(n196), .B2(c[51]), .ZN(n58) );
  INV_X1 U104 ( .A(n59), .ZN(carry[53]) );
  AOI22_X1 U105 ( .A1(b[52]), .A2(a[52]), .B1(n197), .B2(c[52]), .ZN(n59) );
  INV_X1 U106 ( .A(n60), .ZN(carry[54]) );
  AOI22_X1 U107 ( .A1(b[53]), .A2(a[53]), .B1(n198), .B2(c[53]), .ZN(n60) );
  INV_X1 U108 ( .A(n61), .ZN(carry[55]) );
  AOI22_X1 U109 ( .A1(b[54]), .A2(a[54]), .B1(n199), .B2(c[54]), .ZN(n61) );
  INV_X1 U110 ( .A(n62), .ZN(carry[56]) );
  AOI22_X1 U111 ( .A1(b[55]), .A2(a[55]), .B1(n200), .B2(c[55]), .ZN(n62) );
  INV_X1 U112 ( .A(n63), .ZN(carry[57]) );
  AOI22_X1 U113 ( .A1(b[56]), .A2(a[56]), .B1(n201), .B2(c[56]), .ZN(n63) );
  INV_X1 U114 ( .A(n139), .ZN(carry[58]) );
  AOI22_X1 U115 ( .A1(b[57]), .A2(a[57]), .B1(n202), .B2(c[57]), .ZN(n139) );
  INV_X1 U116 ( .A(n140), .ZN(carry[59]) );
  AOI22_X1 U117 ( .A1(b[58]), .A2(a[58]), .B1(n203), .B2(c[58]), .ZN(n140) );
  INV_X1 U118 ( .A(n142), .ZN(carry[60]) );
  AOI22_X1 U119 ( .A1(b[59]), .A2(a[59]), .B1(n204), .B2(c[59]), .ZN(n142) );
  INV_X1 U120 ( .A(n144), .ZN(carry[62]) );
  AOI22_X1 U121 ( .A1(b[61]), .A2(a[61]), .B1(n207), .B2(c[61]), .ZN(n144) );
  INV_X1 U122 ( .A(n145), .ZN(carry[63]) );
  AOI22_X1 U123 ( .A1(b[62]), .A2(a[62]), .B1(n208), .B2(c[62]), .ZN(n145) );
  INV_X1 U124 ( .A(n143), .ZN(carry[61]) );
  AOI22_X1 U125 ( .A1(b[60]), .A2(a[60]), .B1(n206), .B2(c[60]), .ZN(n143) );
  INV_X1 U126 ( .A(n33), .ZN(carry[2]) );
  AOI22_X1 U127 ( .A1(b[1]), .A2(a[1]), .B1(n161), .B2(c[1]), .ZN(n33) );
  INV_X1 U193 ( .A(n44), .ZN(carry[3]) );
  AOI22_X1 U194 ( .A1(b[2]), .A2(a[2]), .B1(n172), .B2(c[2]), .ZN(n44) );
  INV_X1 U195 ( .A(n55), .ZN(carry[4]) );
  AOI22_X1 U253 ( .A1(b[3]), .A2(a[3]), .B1(n183), .B2(c[3]), .ZN(n55) );
  INV_X1 U254 ( .A(n141), .ZN(carry[5]) );
  AOI22_X1 U255 ( .A1(b[4]), .A2(a[4]), .B1(n194), .B2(c[4]), .ZN(n141) );
  INV_X1 U256 ( .A(n146), .ZN(carry[6]) );
  AOI22_X1 U257 ( .A1(b[5]), .A2(a[5]), .B1(n205), .B2(c[5]), .ZN(n146) );
  INV_X1 U258 ( .A(n22), .ZN(carry[1]) );
  AOI22_X1 U259 ( .A1(b[0]), .A2(a[0]), .B1(n150), .B2(c[0]), .ZN(n22) );
  AOI22_X1 U260 ( .A1(b[10]), .A2(a[10]), .B1(n151), .B2(c[10]), .ZN(n13) );
  INV_X1 U261 ( .A(n148), .ZN(carry[8]) );
  AOI22_X1 U262 ( .A1(b[9]), .A2(a[9]), .B1(n213), .B2(c[9]), .ZN(n12) );
  INV_X1 U263 ( .A(n147), .ZN(carry[7]) );
  AOI22_X1 U264 ( .A1(b[6]), .A2(n1), .B1(n210), .B2(c[6]), .ZN(n147) );
  AOI22_X1 U265 ( .A1(b[7]), .A2(n7), .B1(n211), .B2(c[7]), .ZN(n148) );
  AOI22_X1 U266 ( .A1(b[8]), .A2(n2), .B1(n6), .B2(c[8]), .ZN(n149) );
endmodule


module BWAdder_2 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(n211), .B(c[9]), .Z(result[9]) );
  XOR2_X1 U129 ( .A(n210), .B(c[8]), .Z(result[8]) );
  XOR2_X1 U130 ( .A(n209), .B(c[7]), .Z(result[7]) );
  XOR2_X1 U131 ( .A(n208), .B(c[6]), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n207), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n207) );
  XOR2_X1 U134 ( .A(c[62]), .B(n206), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n205), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n204), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n203), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n202), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n201), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n200), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n199), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n198), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n197), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n196), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n195), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n194), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n193), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n192), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n191), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n190), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n189), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n188), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n187), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n186), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n185), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n184), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n183), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n182), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n181), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n180), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n179), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n178), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n177), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n176), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n175), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n174), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n173), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n172), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n171), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n170), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n169), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n168), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n167), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n166), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n165), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n164), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n163), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n162), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n161), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n160), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n159), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n158), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n157), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n156), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n155), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n154), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n153), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n152), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n151), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n150), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n149), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n148), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n210) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n209) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n208) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n203) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n206) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n205) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n204) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n202) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n192) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n201) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n200) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n199) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n198) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n197) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n196) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n195) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n194) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n193) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n191) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n181) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n190) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n189) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n188) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n187) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n186) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n185) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n184) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n183) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n182) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n180) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n170) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n179) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n178) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n177) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n176) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n175) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n174) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n173) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n172) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n171) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n169) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n159) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n168) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n167) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n166) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n165) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n164) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n163) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n162) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n161) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n160) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n158) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n148) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n157) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n156) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n155) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n154) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n153) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n152) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n151) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n150) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n149) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n211) );
  CLKBUF_X1 U2 ( .A(a[10]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(a[5]), .Z(n2) );
  CLKBUF_X1 U4 ( .A(a[9]), .Z(n3) );
  CLKBUF_X1 U5 ( .A(a[8]), .Z(n4) );
  CLKBUF_X1 U6 ( .A(n209), .Z(n5) );
  CLKBUF_X1 U7 ( .A(n149), .Z(n6) );
  CLKBUF_X1 U8 ( .A(n210), .Z(n7) );
  CLKBUF_X1 U9 ( .A(n211), .Z(n8) );
  CLKBUF_X1 U10 ( .A(a[7]), .Z(n9) );
  CLKBUF_X1 U11 ( .A(a[6]), .Z(n10) );
  INV_X1 U12 ( .A(n22), .ZN(carry[20]) );
  AOI22_X1 U13 ( .A1(b[19]), .A2(a[19]), .B1(n158), .B2(c[19]), .ZN(n22) );
  INV_X1 U14 ( .A(n24), .ZN(carry[22]) );
  AOI22_X1 U15 ( .A1(b[21]), .A2(a[21]), .B1(n161), .B2(c[21]), .ZN(n24) );
  INV_X1 U16 ( .A(n26), .ZN(carry[24]) );
  AOI22_X1 U17 ( .A1(b[23]), .A2(a[23]), .B1(n163), .B2(c[23]), .ZN(n26) );
  INV_X1 U18 ( .A(n28), .ZN(carry[26]) );
  AOI22_X1 U19 ( .A1(b[25]), .A2(a[25]), .B1(n165), .B2(c[25]), .ZN(n28) );
  INV_X1 U20 ( .A(n30), .ZN(carry[28]) );
  AOI22_X1 U21 ( .A1(b[27]), .A2(a[27]), .B1(n167), .B2(c[27]), .ZN(n30) );
  INV_X1 U22 ( .A(n33), .ZN(carry[30]) );
  AOI22_X1 U23 ( .A1(b[29]), .A2(a[29]), .B1(n169), .B2(c[29]), .ZN(n33) );
  INV_X1 U24 ( .A(n12), .ZN(carry[11]) );
  INV_X1 U25 ( .A(n23), .ZN(carry[21]) );
  AOI22_X1 U26 ( .A1(b[20]), .A2(a[20]), .B1(n160), .B2(c[20]), .ZN(n23) );
  INV_X1 U27 ( .A(n20), .ZN(carry[19]) );
  AOI22_X1 U28 ( .A1(b[18]), .A2(a[18]), .B1(n157), .B2(c[18]), .ZN(n20) );
  INV_X1 U29 ( .A(n18), .ZN(carry[17]) );
  AOI22_X1 U30 ( .A1(b[16]), .A2(a[16]), .B1(n155), .B2(c[16]), .ZN(n18) );
  INV_X1 U31 ( .A(n19), .ZN(carry[18]) );
  AOI22_X1 U32 ( .A1(b[17]), .A2(a[17]), .B1(n156), .B2(c[17]), .ZN(n19) );
  INV_X1 U33 ( .A(n17), .ZN(carry[16]) );
  AOI22_X1 U34 ( .A1(b[15]), .A2(a[15]), .B1(n154), .B2(c[15]), .ZN(n17) );
  INV_X1 U35 ( .A(n25), .ZN(carry[23]) );
  AOI22_X1 U36 ( .A1(b[22]), .A2(a[22]), .B1(n162), .B2(c[22]), .ZN(n25) );
  INV_X1 U37 ( .A(n27), .ZN(carry[25]) );
  AOI22_X1 U38 ( .A1(b[24]), .A2(a[24]), .B1(n164), .B2(c[24]), .ZN(n27) );
  INV_X1 U39 ( .A(n29), .ZN(carry[27]) );
  AOI22_X1 U40 ( .A1(b[26]), .A2(a[26]), .B1(n166), .B2(c[26]), .ZN(n29) );
  INV_X1 U41 ( .A(n31), .ZN(carry[29]) );
  AOI22_X1 U42 ( .A1(b[28]), .A2(a[28]), .B1(n168), .B2(c[28]), .ZN(n31) );
  INV_X1 U43 ( .A(n34), .ZN(carry[31]) );
  AOI22_X1 U44 ( .A1(b[30]), .A2(a[30]), .B1(n171), .B2(c[30]), .ZN(n34) );
  INV_X1 U45 ( .A(n13), .ZN(carry[12]) );
  AOI22_X1 U46 ( .A1(b[11]), .A2(a[11]), .B1(n150), .B2(c[11]), .ZN(n13) );
  INV_X1 U47 ( .A(n14), .ZN(carry[13]) );
  AOI22_X1 U48 ( .A1(b[12]), .A2(a[12]), .B1(n151), .B2(c[12]), .ZN(n14) );
  INV_X1 U49 ( .A(n15), .ZN(carry[14]) );
  AOI22_X1 U50 ( .A1(b[13]), .A2(a[13]), .B1(n152), .B2(c[13]), .ZN(n15) );
  INV_X1 U51 ( .A(n16), .ZN(carry[15]) );
  AOI22_X1 U52 ( .A1(b[14]), .A2(a[14]), .B1(n153), .B2(c[14]), .ZN(n16) );
  INV_X1 U53 ( .A(n144), .ZN(carry[6]) );
  INV_X1 U54 ( .A(n146), .ZN(carry[8]) );
  INV_X1 U55 ( .A(n145), .ZN(carry[7]) );
  INV_X1 U56 ( .A(n147), .ZN(carry[9]) );
  INV_X1 U57 ( .A(n11), .ZN(carry[10]) );
  INV_X1 U58 ( .A(n35), .ZN(carry[32]) );
  AOI22_X1 U59 ( .A1(b[31]), .A2(a[31]), .B1(n172), .B2(c[31]), .ZN(n35) );
  INV_X1 U60 ( .A(n36), .ZN(carry[33]) );
  AOI22_X1 U61 ( .A1(b[32]), .A2(a[32]), .B1(n173), .B2(c[32]), .ZN(n36) );
  INV_X1 U62 ( .A(n37), .ZN(carry[34]) );
  AOI22_X1 U63 ( .A1(b[33]), .A2(a[33]), .B1(n174), .B2(c[33]), .ZN(n37) );
  INV_X1 U64 ( .A(n39), .ZN(carry[36]) );
  AOI22_X1 U65 ( .A1(b[35]), .A2(a[35]), .B1(n176), .B2(c[35]), .ZN(n39) );
  INV_X1 U66 ( .A(n41), .ZN(carry[38]) );
  AOI22_X1 U67 ( .A1(b[37]), .A2(a[37]), .B1(n178), .B2(c[37]), .ZN(n41) );
  INV_X1 U68 ( .A(n45), .ZN(carry[41]) );
  AOI22_X1 U69 ( .A1(b[40]), .A2(a[40]), .B1(n182), .B2(c[40]), .ZN(n45) );
  INV_X1 U70 ( .A(n46), .ZN(carry[42]) );
  AOI22_X1 U71 ( .A1(b[41]), .A2(a[41]), .B1(n183), .B2(c[41]), .ZN(n46) );
  INV_X1 U72 ( .A(n38), .ZN(carry[35]) );
  AOI22_X1 U73 ( .A1(b[34]), .A2(a[34]), .B1(n175), .B2(c[34]), .ZN(n38) );
  INV_X1 U74 ( .A(n40), .ZN(carry[37]) );
  AOI22_X1 U75 ( .A1(b[36]), .A2(a[36]), .B1(n177), .B2(c[36]), .ZN(n40) );
  INV_X1 U76 ( .A(n42), .ZN(carry[39]) );
  AOI22_X1 U77 ( .A1(b[38]), .A2(a[38]), .B1(n179), .B2(c[38]), .ZN(n42) );
  INV_X1 U78 ( .A(n44), .ZN(carry[40]) );
  AOI22_X1 U79 ( .A1(b[39]), .A2(a[39]), .B1(n180), .B2(c[39]), .ZN(n44) );
  INV_X1 U80 ( .A(n47), .ZN(carry[43]) );
  AOI22_X1 U81 ( .A1(b[42]), .A2(a[42]), .B1(n184), .B2(c[42]), .ZN(n47) );
  INV_X1 U82 ( .A(n48), .ZN(carry[44]) );
  AOI22_X1 U83 ( .A1(b[43]), .A2(a[43]), .B1(n185), .B2(c[43]), .ZN(n48) );
  INV_X1 U84 ( .A(n49), .ZN(carry[45]) );
  AOI22_X1 U85 ( .A1(b[44]), .A2(a[44]), .B1(n186), .B2(c[44]), .ZN(n49) );
  INV_X1 U86 ( .A(n50), .ZN(carry[46]) );
  AOI22_X1 U87 ( .A1(b[45]), .A2(a[45]), .B1(n187), .B2(c[45]), .ZN(n50) );
  INV_X1 U88 ( .A(n51), .ZN(carry[47]) );
  AOI22_X1 U89 ( .A1(b[46]), .A2(a[46]), .B1(n188), .B2(c[46]), .ZN(n51) );
  INV_X1 U90 ( .A(n52), .ZN(carry[48]) );
  AOI22_X1 U91 ( .A1(b[47]), .A2(a[47]), .B1(n189), .B2(c[47]), .ZN(n52) );
  INV_X1 U92 ( .A(n53), .ZN(carry[49]) );
  AOI22_X1 U93 ( .A1(b[48]), .A2(a[48]), .B1(n190), .B2(c[48]), .ZN(n53) );
  INV_X1 U94 ( .A(n55), .ZN(carry[50]) );
  AOI22_X1 U95 ( .A1(b[49]), .A2(a[49]), .B1(n191), .B2(c[49]), .ZN(n55) );
  INV_X1 U96 ( .A(n56), .ZN(carry[51]) );
  AOI22_X1 U97 ( .A1(b[50]), .A2(a[50]), .B1(n193), .B2(c[50]), .ZN(n56) );
  INV_X1 U98 ( .A(n57), .ZN(carry[52]) );
  AOI22_X1 U99 ( .A1(b[51]), .A2(a[51]), .B1(n194), .B2(c[51]), .ZN(n57) );
  INV_X1 U100 ( .A(n58), .ZN(carry[53]) );
  AOI22_X1 U101 ( .A1(b[52]), .A2(a[52]), .B1(n195), .B2(c[52]), .ZN(n58) );
  INV_X1 U102 ( .A(n59), .ZN(carry[54]) );
  AOI22_X1 U103 ( .A1(b[53]), .A2(a[53]), .B1(n196), .B2(c[53]), .ZN(n59) );
  INV_X1 U104 ( .A(n60), .ZN(carry[55]) );
  AOI22_X1 U105 ( .A1(b[54]), .A2(a[54]), .B1(n197), .B2(c[54]), .ZN(n60) );
  INV_X1 U106 ( .A(n61), .ZN(carry[56]) );
  AOI22_X1 U107 ( .A1(b[55]), .A2(a[55]), .B1(n198), .B2(c[55]), .ZN(n61) );
  INV_X1 U108 ( .A(n62), .ZN(carry[57]) );
  AOI22_X1 U109 ( .A1(b[56]), .A2(a[56]), .B1(n199), .B2(c[56]), .ZN(n62) );
  INV_X1 U110 ( .A(n63), .ZN(carry[58]) );
  AOI22_X1 U111 ( .A1(b[57]), .A2(a[57]), .B1(n200), .B2(c[57]), .ZN(n63) );
  INV_X1 U112 ( .A(n138), .ZN(carry[59]) );
  AOI22_X1 U113 ( .A1(b[58]), .A2(a[58]), .B1(n201), .B2(c[58]), .ZN(n138) );
  INV_X1 U114 ( .A(n140), .ZN(carry[60]) );
  AOI22_X1 U115 ( .A1(b[59]), .A2(a[59]), .B1(n202), .B2(c[59]), .ZN(n140) );
  INV_X1 U116 ( .A(n141), .ZN(carry[61]) );
  AOI22_X1 U117 ( .A1(b[60]), .A2(a[60]), .B1(n204), .B2(c[60]), .ZN(n141) );
  INV_X1 U118 ( .A(n142), .ZN(carry[62]) );
  AOI22_X1 U119 ( .A1(b[61]), .A2(a[61]), .B1(n205), .B2(c[61]), .ZN(n142) );
  INV_X1 U120 ( .A(n143), .ZN(carry[63]) );
  AOI22_X1 U121 ( .A1(b[62]), .A2(a[62]), .B1(n206), .B2(c[62]), .ZN(n143) );
  INV_X1 U122 ( .A(n139), .ZN(carry[5]) );
  AOI22_X1 U123 ( .A1(b[4]), .A2(a[4]), .B1(n192), .B2(c[4]), .ZN(n139) );
  INV_X1 U124 ( .A(n54), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n181), .B2(c[3]), .ZN(n54) );
  INV_X1 U126 ( .A(n43), .ZN(carry[3]) );
  AOI22_X1 U127 ( .A1(b[2]), .A2(a[2]), .B1(n170), .B2(c[2]), .ZN(n43) );
  INV_X1 U256 ( .A(n32), .ZN(carry[2]) );
  AOI22_X1 U257 ( .A1(b[1]), .A2(a[1]), .B1(n159), .B2(c[1]), .ZN(n32) );
  INV_X1 U258 ( .A(n21), .ZN(carry[1]) );
  AOI22_X1 U259 ( .A1(b[0]), .A2(a[0]), .B1(n148), .B2(c[0]), .ZN(n21) );
  AOI22_X1 U260 ( .A1(b[6]), .A2(n10), .B1(n208), .B2(c[6]), .ZN(n145) );
  AOI22_X1 U261 ( .A1(b[10]), .A2(n1), .B1(n6), .B2(c[10]), .ZN(n12) );
  AOI22_X1 U262 ( .A1(b[5]), .A2(n2), .B1(n203), .B2(c[5]), .ZN(n144) );
  AOI22_X1 U263 ( .A1(b[9]), .A2(n3), .B1(n8), .B2(c[9]), .ZN(n11) );
  AOI22_X1 U264 ( .A1(b[7]), .A2(n9), .B1(n5), .B2(c[7]), .ZN(n146) );
  AOI22_X1 U265 ( .A1(b[8]), .A2(n4), .B1(n7), .B2(c[8]), .ZN(n147) );
endmodule


module BWAdder_3 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(n201), .B(c[9]), .Z(result[9]) );
  XOR2_X1 U129 ( .A(n200), .B(c[8]), .Z(result[8]) );
  XOR2_X1 U130 ( .A(n199), .B(c[7]), .Z(result[7]) );
  XOR2_X1 U131 ( .A(n198), .B(c[6]), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n197), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n197) );
  XOR2_X1 U134 ( .A(c[62]), .B(n196), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n195), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n194), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n193), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n192), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n191), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n190), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n189), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n188), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n187), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n186), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n185), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n184), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n183), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n182), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n181), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n180), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n179), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n178), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n177), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n176), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n175), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n174), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n173), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n172), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n171), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n170), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n169), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n168), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n167), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n166), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n165), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n164), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n163), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n162), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n161), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n160), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n159), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n158), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n157), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n156), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n155), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n154), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n153), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n152), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n151), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n150), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n149), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n148), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n147), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n146), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n145), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n144), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n143), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n142), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n141), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n140), .Z(result[11]) );
  XOR2_X1 U191 ( .A(n139), .B(c[10]), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n138), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n200) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n199) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n198) );
  XOR2_X1 U196 ( .A(b[5]), .B(a[5]), .Z(n193) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n196) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n195) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n194) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n192) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n182) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n191) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n190) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n189) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n188) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n187) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n186) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n185) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n184) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n183) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n181) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n171) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n180) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n179) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n178) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n177) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n176) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n175) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n174) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n173) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n172) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n170) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n160) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n169) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n168) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n167) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n166) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n165) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n164) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n163) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n162) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n161) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n159) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n149) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n158) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n157) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n156) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n155) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n154) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n153) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n152) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n151) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n150) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n148) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n138) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n147) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n146) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n145) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n144) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n143) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n142) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n141) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n140) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n139) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n201) );
  CLKBUF_X1 U2 ( .A(n199), .Z(n1) );
  CLKBUF_X1 U3 ( .A(b[6]), .Z(n2) );
  CLKBUF_X1 U4 ( .A(n200), .Z(n3) );
  CLKBUF_X1 U5 ( .A(a[8]), .Z(n4) );
  CLKBUF_X1 U6 ( .A(a[6]), .Z(n5) );
  INV_X1 U7 ( .A(n18), .ZN(carry[21]) );
  AOI22_X1 U8 ( .A1(b[20]), .A2(a[20]), .B1(n150), .B2(c[20]), .ZN(n18) );
  INV_X1 U9 ( .A(n17), .ZN(carry[20]) );
  AOI22_X1 U10 ( .A1(b[19]), .A2(a[19]), .B1(n148), .B2(c[19]), .ZN(n17) );
  INV_X1 U11 ( .A(n15), .ZN(carry[19]) );
  AOI22_X1 U12 ( .A1(b[18]), .A2(a[18]), .B1(n147), .B2(c[18]), .ZN(n15) );
  INV_X1 U13 ( .A(n7), .ZN(carry[11]) );
  AOI22_X1 U14 ( .A1(b[10]), .A2(a[10]), .B1(n139), .B2(c[10]), .ZN(n7) );
  INV_X1 U15 ( .A(n8), .ZN(carry[12]) );
  AOI22_X1 U16 ( .A1(b[11]), .A2(a[11]), .B1(n140), .B2(c[11]), .ZN(n8) );
  INV_X1 U17 ( .A(n9), .ZN(carry[13]) );
  AOI22_X1 U18 ( .A1(b[12]), .A2(a[12]), .B1(n141), .B2(c[12]), .ZN(n9) );
  INV_X1 U19 ( .A(n13), .ZN(carry[17]) );
  AOI22_X1 U20 ( .A1(b[16]), .A2(a[16]), .B1(n145), .B2(c[16]), .ZN(n13) );
  INV_X1 U21 ( .A(n10), .ZN(carry[14]) );
  AOI22_X1 U22 ( .A1(b[13]), .A2(a[13]), .B1(n142), .B2(c[13]), .ZN(n10) );
  INV_X1 U23 ( .A(n11), .ZN(carry[15]) );
  AOI22_X1 U24 ( .A1(b[14]), .A2(a[14]), .B1(n143), .B2(c[14]), .ZN(n11) );
  INV_X1 U25 ( .A(n14), .ZN(carry[18]) );
  AOI22_X1 U26 ( .A1(b[17]), .A2(a[17]), .B1(n146), .B2(c[17]), .ZN(n14) );
  INV_X1 U27 ( .A(n12), .ZN(carry[16]) );
  AOI22_X1 U28 ( .A1(b[15]), .A2(a[15]), .B1(n144), .B2(c[15]), .ZN(n12) );
  INV_X1 U29 ( .A(n19), .ZN(carry[22]) );
  AOI22_X1 U30 ( .A1(b[21]), .A2(a[21]), .B1(n151), .B2(c[21]), .ZN(n19) );
  INV_X1 U31 ( .A(n20), .ZN(carry[23]) );
  AOI22_X1 U32 ( .A1(b[22]), .A2(a[22]), .B1(n152), .B2(c[22]), .ZN(n20) );
  INV_X1 U33 ( .A(n21), .ZN(carry[24]) );
  AOI22_X1 U34 ( .A1(b[23]), .A2(a[23]), .B1(n153), .B2(c[23]), .ZN(n21) );
  INV_X1 U35 ( .A(n22), .ZN(carry[25]) );
  AOI22_X1 U36 ( .A1(b[24]), .A2(a[24]), .B1(n154), .B2(c[24]), .ZN(n22) );
  INV_X1 U37 ( .A(n23), .ZN(carry[26]) );
  AOI22_X1 U38 ( .A1(b[25]), .A2(a[25]), .B1(n155), .B2(c[25]), .ZN(n23) );
  INV_X1 U39 ( .A(n24), .ZN(carry[27]) );
  AOI22_X1 U40 ( .A1(b[26]), .A2(a[26]), .B1(n156), .B2(c[26]), .ZN(n24) );
  INV_X1 U41 ( .A(n25), .ZN(carry[28]) );
  AOI22_X1 U42 ( .A1(b[27]), .A2(a[27]), .B1(n157), .B2(c[27]), .ZN(n25) );
  INV_X1 U43 ( .A(n26), .ZN(carry[29]) );
  AOI22_X1 U44 ( .A1(b[28]), .A2(a[28]), .B1(n158), .B2(c[28]), .ZN(n26) );
  INV_X1 U45 ( .A(n28), .ZN(carry[30]) );
  AOI22_X1 U46 ( .A1(b[29]), .A2(a[29]), .B1(n159), .B2(c[29]), .ZN(n28) );
  INV_X1 U47 ( .A(n29), .ZN(carry[31]) );
  AOI22_X1 U48 ( .A1(b[30]), .A2(a[30]), .B1(n161), .B2(c[30]), .ZN(n29) );
  INV_X1 U49 ( .A(n135), .ZN(carry[7]) );
  INV_X1 U50 ( .A(n136), .ZN(carry[8]) );
  INV_X1 U51 ( .A(n137), .ZN(carry[9]) );
  INV_X1 U52 ( .A(n6), .ZN(carry[10]) );
  INV_X1 U53 ( .A(n134), .ZN(carry[6]) );
  INV_X1 U54 ( .A(n60), .ZN(carry[5]) );
  AOI22_X1 U55 ( .A1(b[4]), .A2(a[4]), .B1(n182), .B2(c[4]), .ZN(n60) );
  INV_X1 U56 ( .A(n30), .ZN(carry[32]) );
  AOI22_X1 U57 ( .A1(b[31]), .A2(a[31]), .B1(n162), .B2(c[31]), .ZN(n30) );
  INV_X1 U58 ( .A(n31), .ZN(carry[33]) );
  AOI22_X1 U59 ( .A1(b[32]), .A2(a[32]), .B1(n163), .B2(c[32]), .ZN(n31) );
  INV_X1 U60 ( .A(n32), .ZN(carry[34]) );
  AOI22_X1 U61 ( .A1(b[33]), .A2(a[33]), .B1(n164), .B2(c[33]), .ZN(n32) );
  INV_X1 U62 ( .A(n33), .ZN(carry[35]) );
  AOI22_X1 U63 ( .A1(b[34]), .A2(a[34]), .B1(n165), .B2(c[34]), .ZN(n33) );
  INV_X1 U64 ( .A(n34), .ZN(carry[36]) );
  AOI22_X1 U65 ( .A1(b[35]), .A2(a[35]), .B1(n166), .B2(c[35]), .ZN(n34) );
  INV_X1 U66 ( .A(n35), .ZN(carry[37]) );
  AOI22_X1 U67 ( .A1(b[36]), .A2(a[36]), .B1(n167), .B2(c[36]), .ZN(n35) );
  INV_X1 U68 ( .A(n36), .ZN(carry[38]) );
  AOI22_X1 U69 ( .A1(b[37]), .A2(a[37]), .B1(n168), .B2(c[37]), .ZN(n36) );
  INV_X1 U70 ( .A(n37), .ZN(carry[39]) );
  AOI22_X1 U71 ( .A1(b[38]), .A2(a[38]), .B1(n169), .B2(c[38]), .ZN(n37) );
  INV_X1 U72 ( .A(n39), .ZN(carry[40]) );
  AOI22_X1 U73 ( .A1(b[39]), .A2(a[39]), .B1(n170), .B2(c[39]), .ZN(n39) );
  INV_X1 U74 ( .A(n40), .ZN(carry[41]) );
  AOI22_X1 U75 ( .A1(b[40]), .A2(a[40]), .B1(n172), .B2(c[40]), .ZN(n40) );
  INV_X1 U76 ( .A(n41), .ZN(carry[42]) );
  AOI22_X1 U77 ( .A1(b[41]), .A2(a[41]), .B1(n173), .B2(c[41]), .ZN(n41) );
  INV_X1 U78 ( .A(n42), .ZN(carry[43]) );
  AOI22_X1 U79 ( .A1(b[42]), .A2(a[42]), .B1(n174), .B2(c[42]), .ZN(n42) );
  INV_X1 U80 ( .A(n43), .ZN(carry[44]) );
  AOI22_X1 U81 ( .A1(b[43]), .A2(a[43]), .B1(n175), .B2(c[43]), .ZN(n43) );
  INV_X1 U82 ( .A(n44), .ZN(carry[45]) );
  AOI22_X1 U83 ( .A1(b[44]), .A2(a[44]), .B1(n176), .B2(c[44]), .ZN(n44) );
  INV_X1 U84 ( .A(n45), .ZN(carry[46]) );
  AOI22_X1 U85 ( .A1(b[45]), .A2(a[45]), .B1(n177), .B2(c[45]), .ZN(n45) );
  INV_X1 U86 ( .A(n46), .ZN(carry[47]) );
  AOI22_X1 U87 ( .A1(b[46]), .A2(a[46]), .B1(n178), .B2(c[46]), .ZN(n46) );
  INV_X1 U88 ( .A(n47), .ZN(carry[48]) );
  AOI22_X1 U89 ( .A1(b[47]), .A2(a[47]), .B1(n179), .B2(c[47]), .ZN(n47) );
  INV_X1 U90 ( .A(n48), .ZN(carry[49]) );
  AOI22_X1 U91 ( .A1(b[48]), .A2(a[48]), .B1(n180), .B2(c[48]), .ZN(n48) );
  INV_X1 U92 ( .A(n50), .ZN(carry[50]) );
  AOI22_X1 U93 ( .A1(b[49]), .A2(a[49]), .B1(n181), .B2(c[49]), .ZN(n50) );
  INV_X1 U94 ( .A(n51), .ZN(carry[51]) );
  AOI22_X1 U95 ( .A1(b[50]), .A2(a[50]), .B1(n183), .B2(c[50]), .ZN(n51) );
  INV_X1 U96 ( .A(n52), .ZN(carry[52]) );
  AOI22_X1 U97 ( .A1(b[51]), .A2(a[51]), .B1(n184), .B2(c[51]), .ZN(n52) );
  INV_X1 U98 ( .A(n53), .ZN(carry[53]) );
  AOI22_X1 U99 ( .A1(b[52]), .A2(a[52]), .B1(n185), .B2(c[52]), .ZN(n53) );
  INV_X1 U100 ( .A(n54), .ZN(carry[54]) );
  AOI22_X1 U101 ( .A1(b[53]), .A2(a[53]), .B1(n186), .B2(c[53]), .ZN(n54) );
  INV_X1 U102 ( .A(n55), .ZN(carry[55]) );
  AOI22_X1 U103 ( .A1(b[54]), .A2(a[54]), .B1(n187), .B2(c[54]), .ZN(n55) );
  AOI22_X1 U104 ( .A1(b[62]), .A2(a[62]), .B1(n196), .B2(c[62]), .ZN(n133) );
  INV_X1 U105 ( .A(n56), .ZN(carry[56]) );
  AOI22_X1 U106 ( .A1(b[55]), .A2(a[55]), .B1(n188), .B2(c[55]), .ZN(n56) );
  INV_X1 U107 ( .A(n57), .ZN(carry[57]) );
  AOI22_X1 U108 ( .A1(b[56]), .A2(a[56]), .B1(n189), .B2(c[56]), .ZN(n57) );
  INV_X1 U109 ( .A(n58), .ZN(carry[58]) );
  AOI22_X1 U110 ( .A1(b[57]), .A2(a[57]), .B1(n190), .B2(c[57]), .ZN(n58) );
  INV_X1 U111 ( .A(n59), .ZN(carry[59]) );
  AOI22_X1 U112 ( .A1(b[58]), .A2(a[58]), .B1(n191), .B2(c[58]), .ZN(n59) );
  INV_X1 U113 ( .A(n61), .ZN(carry[60]) );
  AOI22_X1 U114 ( .A1(b[59]), .A2(a[59]), .B1(n192), .B2(c[59]), .ZN(n61) );
  INV_X1 U115 ( .A(n62), .ZN(carry[61]) );
  AOI22_X1 U116 ( .A1(b[60]), .A2(a[60]), .B1(n194), .B2(c[60]), .ZN(n62) );
  INV_X1 U117 ( .A(n63), .ZN(carry[62]) );
  AOI22_X1 U118 ( .A1(b[61]), .A2(a[61]), .B1(n195), .B2(c[61]), .ZN(n63) );
  INV_X1 U119 ( .A(n49), .ZN(carry[4]) );
  AOI22_X1 U120 ( .A1(b[3]), .A2(a[3]), .B1(n171), .B2(c[3]), .ZN(n49) );
  INV_X1 U121 ( .A(n133), .ZN(carry[63]) );
  INV_X1 U122 ( .A(n38), .ZN(carry[3]) );
  AOI22_X1 U123 ( .A1(b[2]), .A2(a[2]), .B1(n160), .B2(c[2]), .ZN(n38) );
  INV_X1 U124 ( .A(n27), .ZN(carry[2]) );
  AOI22_X1 U125 ( .A1(b[1]), .A2(a[1]), .B1(n149), .B2(c[1]), .ZN(n27) );
  INV_X1 U126 ( .A(n16), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n138), .B2(c[0]), .ZN(n16) );
  AOI22_X1 U256 ( .A1(b[9]), .A2(a[9]), .B1(n201), .B2(c[9]), .ZN(n6) );
  AOI22_X1 U257 ( .A1(b[7]), .A2(a[7]), .B1(n1), .B2(c[7]), .ZN(n136) );
  AOI22_X1 U258 ( .A1(b[5]), .A2(a[5]), .B1(n193), .B2(c[5]), .ZN(n134) );
  AOI22_X1 U259 ( .A1(b[8]), .A2(n4), .B1(n3), .B2(c[8]), .ZN(n137) );
  AOI22_X1 U260 ( .A1(n2), .A2(n5), .B1(n198), .B2(c[6]), .ZN(n135) );
endmodule


module BWAdder_4 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207;
  assign carry[0] = 1'b0;

  XOR2_X1 U132 ( .A(a[63]), .B(n203), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n203) );
  XOR2_X1 U134 ( .A(c[62]), .B(n202), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n201), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n200), .Z(result[60]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n198), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n197), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n196), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n195), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n194), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n193), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n192), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n191), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n190), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n189), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n188), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n187), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n186), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n185), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n184), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n183), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n182), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n181), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n180), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n179), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n178), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n177), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n176), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n175), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n174), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n173), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n172), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n171), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n170), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n169), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n168), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n167), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n166), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n165), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n164), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n163), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n162), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n161), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n160), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n159), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n158), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n157), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n156), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n155), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n154), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n153), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n152), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n151), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n150), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n149), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n148), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n147), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n146), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n145), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n144), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n206) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n205) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n204) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n202) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n201) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n200) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n198) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n188) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n197) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n196) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n195) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n194) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n193) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n192) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n191) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n190) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n189) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n187) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n177) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n186) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n185) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n184) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n183) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n182) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n181) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n180) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n179) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n178) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n176) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n166) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n175) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n174) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n173) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n172) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n171) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n170) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n169) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n168) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n167) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n165) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n155) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n164) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n163) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n162) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n161) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n160) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n159) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n158) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n157) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n156) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n154) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n144) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n153) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n152) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n151) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n150) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n149) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n148) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n147) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n146) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n145) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n207) );
  INV_X1 U2 ( .A(b[5]), .ZN(n2) );
  INV_X1 U3 ( .A(c[9]), .ZN(n3) );
  INV_X1 U4 ( .A(c[7]), .ZN(n7) );
  INV_X1 U5 ( .A(c[6]), .ZN(n6) );
  INV_X1 U6 ( .A(c[5]), .ZN(n5) );
  CLKBUF_X1 U7 ( .A(n205), .Z(n1) );
  XNOR2_X1 U8 ( .A(a[5]), .B(n2), .ZN(n199) );
  XNOR2_X1 U9 ( .A(n3), .B(n207), .ZN(result[9]) );
  CLKBUF_X1 U10 ( .A(a[5]), .Z(n4) );
  XNOR2_X1 U11 ( .A(n5), .B(n199), .ZN(result[5]) );
  XNOR2_X1 U12 ( .A(n204), .B(n6), .ZN(result[6]) );
  XNOR2_X1 U13 ( .A(n205), .B(n7), .ZN(result[7]) );
  XOR2_X1 U14 ( .A(c[8]), .B(n206), .Z(result[8]) );
  INV_X1 U15 ( .A(n16), .ZN(carry[17]) );
  AOI22_X1 U16 ( .A1(b[16]), .A2(a[16]), .B1(n151), .B2(c[16]), .ZN(n16) );
  INV_X1 U17 ( .A(n17), .ZN(carry[18]) );
  AOI22_X1 U18 ( .A1(b[17]), .A2(a[17]), .B1(n152), .B2(c[17]), .ZN(n17) );
  INV_X1 U19 ( .A(n18), .ZN(carry[19]) );
  AOI22_X1 U20 ( .A1(b[18]), .A2(a[18]), .B1(n153), .B2(c[18]), .ZN(n18) );
  INV_X1 U21 ( .A(n20), .ZN(carry[20]) );
  AOI22_X1 U22 ( .A1(b[19]), .A2(a[19]), .B1(n154), .B2(c[19]), .ZN(n20) );
  INV_X1 U23 ( .A(n21), .ZN(carry[21]) );
  AOI22_X1 U24 ( .A1(b[20]), .A2(a[20]), .B1(n156), .B2(c[20]), .ZN(n21) );
  INV_X1 U25 ( .A(n22), .ZN(carry[22]) );
  AOI22_X1 U26 ( .A1(b[21]), .A2(a[21]), .B1(n157), .B2(c[21]), .ZN(n22) );
  INV_X1 U27 ( .A(n23), .ZN(carry[23]) );
  AOI22_X1 U28 ( .A1(b[22]), .A2(a[22]), .B1(n158), .B2(c[22]), .ZN(n23) );
  INV_X1 U29 ( .A(n24), .ZN(carry[24]) );
  AOI22_X1 U30 ( .A1(b[23]), .A2(a[23]), .B1(n159), .B2(c[23]), .ZN(n24) );
  INV_X1 U31 ( .A(n25), .ZN(carry[25]) );
  AOI22_X1 U32 ( .A1(b[24]), .A2(a[24]), .B1(n160), .B2(c[24]), .ZN(n25) );
  INV_X1 U33 ( .A(n26), .ZN(carry[26]) );
  AOI22_X1 U34 ( .A1(b[25]), .A2(a[25]), .B1(n161), .B2(c[25]), .ZN(n26) );
  INV_X1 U35 ( .A(n27), .ZN(carry[27]) );
  AOI22_X1 U36 ( .A1(b[26]), .A2(a[26]), .B1(n162), .B2(c[26]), .ZN(n27) );
  INV_X1 U37 ( .A(n28), .ZN(carry[28]) );
  AOI22_X1 U38 ( .A1(b[27]), .A2(a[27]), .B1(n163), .B2(c[27]), .ZN(n28) );
  INV_X1 U39 ( .A(n29), .ZN(carry[29]) );
  AOI22_X1 U40 ( .A1(b[28]), .A2(a[28]), .B1(n164), .B2(c[28]), .ZN(n29) );
  INV_X1 U41 ( .A(n15), .ZN(carry[16]) );
  AOI22_X1 U42 ( .A1(b[15]), .A2(a[15]), .B1(n150), .B2(c[15]), .ZN(n15) );
  INV_X1 U43 ( .A(n14), .ZN(carry[15]) );
  AOI22_X1 U44 ( .A1(b[14]), .A2(a[14]), .B1(n149), .B2(c[14]), .ZN(n14) );
  INV_X1 U45 ( .A(n35), .ZN(carry[34]) );
  AOI22_X1 U46 ( .A1(b[33]), .A2(a[33]), .B1(n170), .B2(c[33]), .ZN(n35) );
  INV_X1 U47 ( .A(n36), .ZN(carry[35]) );
  AOI22_X1 U48 ( .A1(b[34]), .A2(a[34]), .B1(n171), .B2(c[34]), .ZN(n36) );
  INV_X1 U49 ( .A(n37), .ZN(carry[36]) );
  AOI22_X1 U50 ( .A1(b[35]), .A2(a[35]), .B1(n172), .B2(c[35]), .ZN(n37) );
  INV_X1 U51 ( .A(n38), .ZN(carry[37]) );
  AOI22_X1 U52 ( .A1(b[36]), .A2(a[36]), .B1(n173), .B2(c[36]), .ZN(n38) );
  INV_X1 U53 ( .A(n39), .ZN(carry[38]) );
  AOI22_X1 U54 ( .A1(b[37]), .A2(a[37]), .B1(n174), .B2(c[37]), .ZN(n39) );
  INV_X1 U55 ( .A(n40), .ZN(carry[39]) );
  AOI22_X1 U56 ( .A1(b[38]), .A2(a[38]), .B1(n175), .B2(c[38]), .ZN(n40) );
  INV_X1 U57 ( .A(n42), .ZN(carry[40]) );
  AOI22_X1 U58 ( .A1(b[39]), .A2(a[39]), .B1(n176), .B2(c[39]), .ZN(n42) );
  INV_X1 U59 ( .A(n43), .ZN(carry[41]) );
  AOI22_X1 U60 ( .A1(b[40]), .A2(a[40]), .B1(n178), .B2(c[40]), .ZN(n43) );
  INV_X1 U61 ( .A(n44), .ZN(carry[42]) );
  AOI22_X1 U62 ( .A1(b[41]), .A2(a[41]), .B1(n179), .B2(c[41]), .ZN(n44) );
  INV_X1 U63 ( .A(n34), .ZN(carry[33]) );
  AOI22_X1 U64 ( .A1(b[32]), .A2(a[32]), .B1(n169), .B2(c[32]), .ZN(n34) );
  INV_X1 U65 ( .A(n31), .ZN(carry[30]) );
  AOI22_X1 U66 ( .A1(b[29]), .A2(a[29]), .B1(n165), .B2(c[29]), .ZN(n31) );
  INV_X1 U67 ( .A(n32), .ZN(carry[31]) );
  AOI22_X1 U68 ( .A1(b[30]), .A2(a[30]), .B1(n167), .B2(c[30]), .ZN(n32) );
  INV_X1 U69 ( .A(n33), .ZN(carry[32]) );
  AOI22_X1 U70 ( .A1(b[31]), .A2(a[31]), .B1(n168), .B2(c[31]), .ZN(n33) );
  INV_X1 U71 ( .A(n45), .ZN(carry[43]) );
  AOI22_X1 U72 ( .A1(b[42]), .A2(a[42]), .B1(n180), .B2(c[42]), .ZN(n45) );
  INV_X1 U73 ( .A(n47), .ZN(carry[45]) );
  AOI22_X1 U74 ( .A1(b[44]), .A2(a[44]), .B1(n182), .B2(c[44]), .ZN(n47) );
  INV_X1 U75 ( .A(n50), .ZN(carry[48]) );
  AOI22_X1 U76 ( .A1(b[47]), .A2(a[47]), .B1(n185), .B2(c[47]), .ZN(n50) );
  INV_X1 U77 ( .A(n46), .ZN(carry[44]) );
  AOI22_X1 U78 ( .A1(b[43]), .A2(a[43]), .B1(n181), .B2(c[43]), .ZN(n46) );
  INV_X1 U79 ( .A(n48), .ZN(carry[46]) );
  AOI22_X1 U80 ( .A1(b[45]), .A2(a[45]), .B1(n183), .B2(c[45]), .ZN(n48) );
  INV_X1 U81 ( .A(n49), .ZN(carry[47]) );
  AOI22_X1 U82 ( .A1(b[46]), .A2(a[46]), .B1(n184), .B2(c[46]), .ZN(n49) );
  INV_X1 U83 ( .A(n51), .ZN(carry[49]) );
  AOI22_X1 U84 ( .A1(b[48]), .A2(a[48]), .B1(n186), .B2(c[48]), .ZN(n51) );
  INV_X1 U85 ( .A(n53), .ZN(carry[50]) );
  AOI22_X1 U86 ( .A1(b[49]), .A2(a[49]), .B1(n187), .B2(c[49]), .ZN(n53) );
  INV_X1 U87 ( .A(n54), .ZN(carry[51]) );
  AOI22_X1 U88 ( .A1(b[50]), .A2(a[50]), .B1(n189), .B2(c[50]), .ZN(n54) );
  INV_X1 U89 ( .A(n55), .ZN(carry[52]) );
  AOI22_X1 U90 ( .A1(b[51]), .A2(a[51]), .B1(n190), .B2(c[51]), .ZN(n55) );
  INV_X1 U91 ( .A(n56), .ZN(carry[53]) );
  AOI22_X1 U92 ( .A1(b[52]), .A2(a[52]), .B1(n191), .B2(c[52]), .ZN(n56) );
  INV_X1 U93 ( .A(n57), .ZN(carry[54]) );
  AOI22_X1 U94 ( .A1(b[53]), .A2(a[53]), .B1(n192), .B2(c[53]), .ZN(n57) );
  INV_X1 U95 ( .A(n58), .ZN(carry[55]) );
  AOI22_X1 U96 ( .A1(b[54]), .A2(a[54]), .B1(n193), .B2(c[54]), .ZN(n58) );
  INV_X1 U97 ( .A(n59), .ZN(carry[56]) );
  AOI22_X1 U98 ( .A1(b[55]), .A2(a[55]), .B1(n194), .B2(c[55]), .ZN(n59) );
  INV_X1 U99 ( .A(n60), .ZN(carry[57]) );
  AOI22_X1 U100 ( .A1(b[56]), .A2(a[56]), .B1(n195), .B2(c[56]), .ZN(n60) );
  INV_X1 U101 ( .A(n61), .ZN(carry[58]) );
  AOI22_X1 U102 ( .A1(b[57]), .A2(a[57]), .B1(n196), .B2(c[57]), .ZN(n61) );
  INV_X1 U103 ( .A(n62), .ZN(carry[59]) );
  AOI22_X1 U104 ( .A1(b[58]), .A2(a[58]), .B1(n197), .B2(c[58]), .ZN(n62) );
  INV_X1 U105 ( .A(n136), .ZN(carry[60]) );
  AOI22_X1 U106 ( .A1(b[59]), .A2(a[59]), .B1(n198), .B2(c[59]), .ZN(n136) );
  INV_X1 U107 ( .A(n137), .ZN(carry[61]) );
  AOI22_X1 U108 ( .A1(b[60]), .A2(a[60]), .B1(n200), .B2(c[60]), .ZN(n137) );
  INV_X1 U109 ( .A(n138), .ZN(carry[62]) );
  AOI22_X1 U110 ( .A1(b[61]), .A2(a[61]), .B1(n201), .B2(c[61]), .ZN(n138) );
  INV_X1 U111 ( .A(n139), .ZN(carry[63]) );
  AOI22_X1 U112 ( .A1(b[62]), .A2(a[62]), .B1(n202), .B2(c[62]), .ZN(n139) );
  INV_X1 U113 ( .A(n10), .ZN(carry[11]) );
  AOI22_X1 U114 ( .A1(b[10]), .A2(a[10]), .B1(n145), .B2(c[10]), .ZN(n10) );
  INV_X1 U115 ( .A(n11), .ZN(carry[12]) );
  AOI22_X1 U116 ( .A1(b[11]), .A2(a[11]), .B1(n146), .B2(c[11]), .ZN(n11) );
  INV_X1 U117 ( .A(n12), .ZN(carry[13]) );
  AOI22_X1 U118 ( .A1(b[12]), .A2(a[12]), .B1(n147), .B2(c[12]), .ZN(n12) );
  INV_X1 U119 ( .A(n13), .ZN(carry[14]) );
  AOI22_X1 U120 ( .A1(b[13]), .A2(a[13]), .B1(n148), .B2(c[13]), .ZN(n13) );
  INV_X1 U121 ( .A(n52), .ZN(carry[4]) );
  AOI22_X1 U122 ( .A1(b[3]), .A2(a[3]), .B1(n177), .B2(c[3]), .ZN(n52) );
  INV_X1 U123 ( .A(n140), .ZN(carry[6]) );
  INV_X1 U124 ( .A(n141), .ZN(carry[7]) );
  INV_X1 U125 ( .A(n142), .ZN(carry[8]) );
  INV_X1 U126 ( .A(n143), .ZN(carry[9]) );
  AOI22_X1 U127 ( .A1(b[8]), .A2(a[8]), .B1(n206), .B2(c[8]), .ZN(n143) );
  INV_X1 U128 ( .A(n63), .ZN(carry[5]) );
  AOI22_X1 U129 ( .A1(b[4]), .A2(a[4]), .B1(n188), .B2(c[4]), .ZN(n63) );
  INV_X1 U130 ( .A(n9), .ZN(carry[10]) );
  AOI22_X1 U131 ( .A1(b[9]), .A2(a[9]), .B1(n207), .B2(c[9]), .ZN(n9) );
  INV_X1 U137 ( .A(n41), .ZN(carry[3]) );
  AOI22_X1 U196 ( .A1(b[2]), .A2(a[2]), .B1(n166), .B2(c[2]), .ZN(n41) );
  INV_X1 U256 ( .A(n30), .ZN(carry[2]) );
  AOI22_X1 U257 ( .A1(b[1]), .A2(a[1]), .B1(n155), .B2(c[1]), .ZN(n30) );
  INV_X1 U258 ( .A(n19), .ZN(carry[1]) );
  AOI22_X1 U259 ( .A1(b[0]), .A2(a[0]), .B1(n144), .B2(c[0]), .ZN(n19) );
  CLKBUF_X1 U260 ( .A(a[6]), .Z(n8) );
  AOI22_X1 U261 ( .A1(b[6]), .A2(n8), .B1(n204), .B2(c[6]), .ZN(n141) );
  AOI22_X1 U262 ( .A1(b[5]), .A2(n4), .B1(n199), .B2(c[5]), .ZN(n140) );
  AOI22_X1 U263 ( .A1(b[7]), .A2(a[7]), .B1(n1), .B2(c[7]), .ZN(n142) );
endmodule


module BWAdder_5 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219;
  assign carry[0] = 1'b0;

  XOR2_X1 U132 ( .A(a[63]), .B(n215), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n215) );
  XOR2_X1 U134 ( .A(c[62]), .B(n214), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n213), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n212), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n211), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n210), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n209), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n208), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n207), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n206), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n205), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n204), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n203), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n202), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n201), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n200), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n199), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n198), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n197), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n196), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n195), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n194), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n193), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n192), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n191), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n190), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n189), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n188), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n187), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n186), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n185), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n184), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n183), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n182), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n181), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n180), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n179), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n178), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n177), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n176), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n175), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n174), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n173), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n172), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n171), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n170), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n169), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n168), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n167), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n166), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n165), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n164), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n163), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n162), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n161), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n160), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n159), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n158), .Z(result[11]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n156), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n218) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n217) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n216) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n211) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n214) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n213) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n212) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n210) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n200) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n209) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n208) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n207) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n206) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n205) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n204) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n203) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n202) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n201) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n199) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n189) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n198) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n197) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n196) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n195) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n194) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n193) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n192) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n191) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n190) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n188) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n178) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n187) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n186) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n185) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n184) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n183) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n182) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n181) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n180) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n179) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n177) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n167) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n176) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n175) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n174) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n173) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n172) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n171) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n170) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n169) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n168) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n166) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n156) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n165) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n164) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n163) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n162) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n161) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n160) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n159) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n158) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n157) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n219) );
  CLKBUF_X1 U2 ( .A(n217), .Z(n1) );
  CLKBUF_X1 U3 ( .A(b[8]), .Z(n2) );
  CLKBUF_X1 U4 ( .A(n218), .Z(n3) );
  CLKBUF_X1 U5 ( .A(a[7]), .Z(n4) );
  INV_X1 U6 ( .A(c[10]), .ZN(n6) );
  INV_X1 U7 ( .A(c[6]), .ZN(n7) );
  INV_X1 U8 ( .A(c[7]), .ZN(n8) );
  INV_X1 U9 ( .A(c[8]), .ZN(n14) );
  INV_X1 U10 ( .A(c[9]), .ZN(n12) );
  CLKBUF_X1 U11 ( .A(b[7]), .Z(n5) );
  XNOR2_X1 U12 ( .A(n157), .B(n6), .ZN(result[10]) );
  XNOR2_X1 U13 ( .A(n216), .B(n7), .ZN(result[6]) );
  XNOR2_X1 U14 ( .A(n217), .B(n8), .ZN(result[7]) );
  CLKBUF_X1 U15 ( .A(a[8]), .Z(n9) );
  CLKBUF_X1 U16 ( .A(a[10]), .Z(n10) );
  CLKBUF_X1 U17 ( .A(a[6]), .Z(n11) );
  XNOR2_X1 U18 ( .A(n219), .B(n12), .ZN(result[9]) );
  CLKBUF_X1 U19 ( .A(n216), .Z(n13) );
  XNOR2_X1 U20 ( .A(n218), .B(n14), .ZN(result[8]) );
  INV_X1 U21 ( .A(n151), .ZN(carry[63]) );
  INV_X1 U22 ( .A(n16), .ZN(carry[11]) );
  INV_X1 U23 ( .A(n15), .ZN(carry[10]) );
  INV_X1 U24 ( .A(n29), .ZN(carry[23]) );
  AOI22_X1 U25 ( .A1(b[22]), .A2(a[22]), .B1(n170), .B2(c[22]), .ZN(n29) );
  INV_X1 U26 ( .A(n30), .ZN(carry[24]) );
  AOI22_X1 U27 ( .A1(b[23]), .A2(a[23]), .B1(n171), .B2(c[23]), .ZN(n30) );
  INV_X1 U28 ( .A(n31), .ZN(carry[25]) );
  AOI22_X1 U29 ( .A1(b[24]), .A2(a[24]), .B1(n172), .B2(c[24]), .ZN(n31) );
  INV_X1 U30 ( .A(n32), .ZN(carry[26]) );
  AOI22_X1 U31 ( .A1(b[25]), .A2(a[25]), .B1(n173), .B2(c[25]), .ZN(n32) );
  INV_X1 U32 ( .A(n33), .ZN(carry[27]) );
  AOI22_X1 U33 ( .A1(b[26]), .A2(a[26]), .B1(n174), .B2(c[26]), .ZN(n33) );
  INV_X1 U34 ( .A(n34), .ZN(carry[28]) );
  AOI22_X1 U35 ( .A1(b[27]), .A2(a[27]), .B1(n175), .B2(c[27]), .ZN(n34) );
  INV_X1 U36 ( .A(n35), .ZN(carry[29]) );
  AOI22_X1 U37 ( .A1(b[28]), .A2(a[28]), .B1(n176), .B2(c[28]), .ZN(n35) );
  INV_X1 U38 ( .A(n37), .ZN(carry[30]) );
  AOI22_X1 U39 ( .A1(b[29]), .A2(a[29]), .B1(n177), .B2(c[29]), .ZN(n37) );
  INV_X1 U40 ( .A(n38), .ZN(carry[31]) );
  AOI22_X1 U41 ( .A1(b[30]), .A2(a[30]), .B1(n179), .B2(c[30]), .ZN(n38) );
  INV_X1 U42 ( .A(n26), .ZN(carry[20]) );
  AOI22_X1 U43 ( .A1(b[19]), .A2(a[19]), .B1(n166), .B2(c[19]), .ZN(n26) );
  INV_X1 U44 ( .A(n24), .ZN(carry[19]) );
  AOI22_X1 U45 ( .A1(b[18]), .A2(a[18]), .B1(n165), .B2(c[18]), .ZN(n24) );
  INV_X1 U46 ( .A(n23), .ZN(carry[18]) );
  AOI22_X1 U47 ( .A1(b[17]), .A2(a[17]), .B1(n164), .B2(c[17]), .ZN(n23) );
  INV_X1 U48 ( .A(n22), .ZN(carry[17]) );
  AOI22_X1 U49 ( .A1(b[16]), .A2(a[16]), .B1(n163), .B2(c[16]), .ZN(n22) );
  INV_X1 U50 ( .A(n21), .ZN(carry[16]) );
  AOI22_X1 U51 ( .A1(b[15]), .A2(a[15]), .B1(n162), .B2(c[15]), .ZN(n21) );
  INV_X1 U52 ( .A(n27), .ZN(carry[21]) );
  AOI22_X1 U53 ( .A1(b[20]), .A2(a[20]), .B1(n168), .B2(c[20]), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(carry[22]) );
  AOI22_X1 U55 ( .A1(b[21]), .A2(a[21]), .B1(n169), .B2(c[21]), .ZN(n28) );
  INV_X1 U56 ( .A(n17), .ZN(carry[12]) );
  AOI22_X1 U57 ( .A1(b[11]), .A2(a[11]), .B1(n158), .B2(c[11]), .ZN(n17) );
  INV_X1 U58 ( .A(n18), .ZN(carry[13]) );
  AOI22_X1 U59 ( .A1(b[12]), .A2(a[12]), .B1(n159), .B2(c[12]), .ZN(n18) );
  INV_X1 U60 ( .A(n19), .ZN(carry[14]) );
  AOI22_X1 U61 ( .A1(b[13]), .A2(a[13]), .B1(n160), .B2(c[13]), .ZN(n19) );
  INV_X1 U62 ( .A(n20), .ZN(carry[15]) );
  AOI22_X1 U63 ( .A1(b[14]), .A2(a[14]), .B1(n161), .B2(c[14]), .ZN(n20) );
  INV_X1 U64 ( .A(n153), .ZN(carry[7]) );
  INV_X1 U65 ( .A(n154), .ZN(carry[8]) );
  INV_X1 U66 ( .A(n155), .ZN(carry[9]) );
  INV_X1 U67 ( .A(n152), .ZN(carry[6]) );
  AOI22_X1 U68 ( .A1(b[5]), .A2(a[5]), .B1(n211), .B2(c[5]), .ZN(n152) );
  INV_X1 U69 ( .A(n39), .ZN(carry[32]) );
  AOI22_X1 U70 ( .A1(b[31]), .A2(a[31]), .B1(n180), .B2(c[31]), .ZN(n39) );
  INV_X1 U71 ( .A(n40), .ZN(carry[33]) );
  AOI22_X1 U72 ( .A1(b[32]), .A2(a[32]), .B1(n181), .B2(c[32]), .ZN(n40) );
  INV_X1 U73 ( .A(n41), .ZN(carry[34]) );
  AOI22_X1 U74 ( .A1(b[33]), .A2(a[33]), .B1(n182), .B2(c[33]), .ZN(n41) );
  INV_X1 U75 ( .A(n42), .ZN(carry[35]) );
  AOI22_X1 U76 ( .A1(b[34]), .A2(a[34]), .B1(n183), .B2(c[34]), .ZN(n42) );
  INV_X1 U77 ( .A(n43), .ZN(carry[36]) );
  AOI22_X1 U78 ( .A1(b[35]), .A2(a[35]), .B1(n184), .B2(c[35]), .ZN(n43) );
  INV_X1 U79 ( .A(n44), .ZN(carry[37]) );
  AOI22_X1 U80 ( .A1(b[36]), .A2(a[36]), .B1(n185), .B2(c[36]), .ZN(n44) );
  INV_X1 U81 ( .A(n45), .ZN(carry[38]) );
  AOI22_X1 U82 ( .A1(b[37]), .A2(a[37]), .B1(n186), .B2(c[37]), .ZN(n45) );
  INV_X1 U83 ( .A(n46), .ZN(carry[39]) );
  AOI22_X1 U84 ( .A1(b[38]), .A2(a[38]), .B1(n187), .B2(c[38]), .ZN(n46) );
  INV_X1 U85 ( .A(n48), .ZN(carry[40]) );
  AOI22_X1 U86 ( .A1(b[39]), .A2(a[39]), .B1(n188), .B2(c[39]), .ZN(n48) );
  INV_X1 U87 ( .A(n49), .ZN(carry[41]) );
  AOI22_X1 U88 ( .A1(b[40]), .A2(a[40]), .B1(n190), .B2(c[40]), .ZN(n49) );
  INV_X1 U89 ( .A(n50), .ZN(carry[42]) );
  AOI22_X1 U90 ( .A1(b[41]), .A2(a[41]), .B1(n191), .B2(c[41]), .ZN(n50) );
  INV_X1 U91 ( .A(n51), .ZN(carry[43]) );
  AOI22_X1 U92 ( .A1(b[42]), .A2(a[42]), .B1(n192), .B2(c[42]), .ZN(n51) );
  INV_X1 U93 ( .A(n52), .ZN(carry[44]) );
  AOI22_X1 U94 ( .A1(b[43]), .A2(a[43]), .B1(n193), .B2(c[43]), .ZN(n52) );
  INV_X1 U95 ( .A(n53), .ZN(carry[45]) );
  AOI22_X1 U96 ( .A1(b[44]), .A2(a[44]), .B1(n194), .B2(c[44]), .ZN(n53) );
  INV_X1 U97 ( .A(n54), .ZN(carry[46]) );
  AOI22_X1 U98 ( .A1(b[45]), .A2(a[45]), .B1(n195), .B2(c[45]), .ZN(n54) );
  INV_X1 U99 ( .A(n55), .ZN(carry[47]) );
  AOI22_X1 U100 ( .A1(b[46]), .A2(a[46]), .B1(n196), .B2(c[46]), .ZN(n55) );
  INV_X1 U101 ( .A(n56), .ZN(carry[48]) );
  AOI22_X1 U102 ( .A1(b[47]), .A2(a[47]), .B1(n197), .B2(c[47]), .ZN(n56) );
  INV_X1 U103 ( .A(n57), .ZN(carry[49]) );
  AOI22_X1 U104 ( .A1(b[48]), .A2(a[48]), .B1(n198), .B2(c[48]), .ZN(n57) );
  INV_X1 U105 ( .A(n59), .ZN(carry[50]) );
  AOI22_X1 U106 ( .A1(b[49]), .A2(a[49]), .B1(n199), .B2(c[49]), .ZN(n59) );
  INV_X1 U107 ( .A(n60), .ZN(carry[51]) );
  AOI22_X1 U108 ( .A1(b[50]), .A2(a[50]), .B1(n201), .B2(c[50]), .ZN(n60) );
  INV_X1 U109 ( .A(n61), .ZN(carry[52]) );
  AOI22_X1 U110 ( .A1(b[51]), .A2(a[51]), .B1(n202), .B2(c[51]), .ZN(n61) );
  INV_X1 U111 ( .A(n62), .ZN(carry[53]) );
  AOI22_X1 U112 ( .A1(b[52]), .A2(a[52]), .B1(n203), .B2(c[52]), .ZN(n62) );
  INV_X1 U113 ( .A(n63), .ZN(carry[54]) );
  AOI22_X1 U114 ( .A1(b[53]), .A2(a[53]), .B1(n204), .B2(c[53]), .ZN(n63) );
  INV_X1 U115 ( .A(n142), .ZN(carry[55]) );
  AOI22_X1 U116 ( .A1(b[54]), .A2(a[54]), .B1(n205), .B2(c[54]), .ZN(n142) );
  AOI22_X1 U117 ( .A1(b[62]), .A2(a[62]), .B1(n214), .B2(c[62]), .ZN(n151) );
  INV_X1 U118 ( .A(n143), .ZN(carry[56]) );
  AOI22_X1 U119 ( .A1(b[55]), .A2(a[55]), .B1(n206), .B2(c[55]), .ZN(n143) );
  INV_X1 U120 ( .A(n144), .ZN(carry[57]) );
  AOI22_X1 U121 ( .A1(b[56]), .A2(a[56]), .B1(n207), .B2(c[56]), .ZN(n144) );
  INV_X1 U122 ( .A(n145), .ZN(carry[58]) );
  AOI22_X1 U123 ( .A1(b[57]), .A2(a[57]), .B1(n208), .B2(c[57]), .ZN(n145) );
  INV_X1 U124 ( .A(n146), .ZN(carry[59]) );
  AOI22_X1 U125 ( .A1(b[58]), .A2(a[58]), .B1(n209), .B2(c[58]), .ZN(n146) );
  INV_X1 U126 ( .A(n148), .ZN(carry[60]) );
  AOI22_X1 U127 ( .A1(b[59]), .A2(a[59]), .B1(n210), .B2(c[59]), .ZN(n148) );
  INV_X1 U128 ( .A(n149), .ZN(carry[61]) );
  AOI22_X1 U129 ( .A1(b[60]), .A2(a[60]), .B1(n212), .B2(c[60]), .ZN(n149) );
  INV_X1 U130 ( .A(n150), .ZN(carry[62]) );
  AOI22_X1 U131 ( .A1(b[61]), .A2(a[61]), .B1(n213), .B2(c[61]), .ZN(n150) );
  INV_X1 U191 ( .A(n47), .ZN(carry[3]) );
  AOI22_X1 U256 ( .A1(b[2]), .A2(a[2]), .B1(n178), .B2(c[2]), .ZN(n47) );
  INV_X1 U257 ( .A(n58), .ZN(carry[4]) );
  AOI22_X1 U258 ( .A1(b[3]), .A2(a[3]), .B1(n189), .B2(c[3]), .ZN(n58) );
  INV_X1 U259 ( .A(n147), .ZN(carry[5]) );
  AOI22_X1 U260 ( .A1(b[4]), .A2(a[4]), .B1(n200), .B2(c[4]), .ZN(n147) );
  INV_X1 U261 ( .A(n36), .ZN(carry[2]) );
  AOI22_X1 U262 ( .A1(b[1]), .A2(a[1]), .B1(n167), .B2(c[1]), .ZN(n36) );
  INV_X1 U263 ( .A(n25), .ZN(carry[1]) );
  AOI22_X1 U264 ( .A1(b[0]), .A2(a[0]), .B1(n156), .B2(c[0]), .ZN(n25) );
  AOI22_X1 U265 ( .A1(b[10]), .A2(n10), .B1(n157), .B2(c[10]), .ZN(n16) );
  AOI22_X1 U266 ( .A1(b[9]), .A2(a[9]), .B1(n219), .B2(c[9]), .ZN(n15) );
  AOI22_X1 U267 ( .A1(b[6]), .A2(n11), .B1(n13), .B2(c[6]), .ZN(n153) );
  AOI22_X1 U268 ( .A1(n2), .A2(n9), .B1(n3), .B2(c[8]), .ZN(n155) );
  AOI22_X1 U269 ( .A1(n5), .A2(n4), .B1(n1), .B2(c[7]), .ZN(n154) );
endmodule


module BWAdder_6 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n59), .ZN(carry[63]) );
  INV_X1 U3 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U4 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U5 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U6 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U7 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U8 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U9 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U10 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U11 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U12 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U13 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U14 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U15 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U16 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U17 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U18 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U19 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U20 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U21 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U22 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U23 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U24 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U25 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U26 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U27 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U28 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U29 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U30 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U31 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U32 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U33 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U34 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U35 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U36 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U37 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U38 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U39 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U40 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U41 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U42 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U43 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U44 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U45 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U46 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  AOI22_X1 U47 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U48 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U49 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U50 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U51 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U52 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U53 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U54 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U55 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U56 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U57 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U58 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U59 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U60 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U61 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U62 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U63 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U64 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U65 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U66 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U67 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U68 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U69 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U70 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U71 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U72 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U73 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U74 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U75 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U76 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U77 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U78 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U79 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U80 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U81 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U82 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U83 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U84 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U85 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U86 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U87 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U88 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U89 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U90 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U91 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U92 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U93 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U94 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U95 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U96 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U97 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U98 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U99 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U100 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U101 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U102 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U103 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U104 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U105 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U106 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U107 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U108 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U109 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U110 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U111 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U112 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U113 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U114 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U115 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U116 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U117 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U118 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U119 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U120 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U121 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U122 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U123 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U124 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U125 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_7 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n199), .Z(result[9]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n196), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n195), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n195) );
  XOR2_X1 U134 ( .A(c[62]), .B(n194), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n193), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n192), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n191), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n190), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n189), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n188), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n187), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n186), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n185), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n184), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n183), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n182), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n181), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n180), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n179), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n178), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n177), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n176), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n175), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n174), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n173), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n172), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n171), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n170), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n169), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n168), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n167), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n166), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n165), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n164), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n163), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n162), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n161), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n160), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n159), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n158), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n157), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n156), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n155), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n154), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n153), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n152), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n151), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n150), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n149), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n148), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n147), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n146), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n145), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n144), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n143), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n142), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n141), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n140), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n139), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n138), .Z(result[11]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n136), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n198) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n196) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n191) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n194) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n193) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n192) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n190) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n180) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n189) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n188) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n187) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n186) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n185) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n184) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n183) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n182) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n181) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n179) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n169) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n178) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n177) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n176) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n175) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n174) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n173) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n172) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n171) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n170) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n168) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n158) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n167) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n166) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n165) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n164) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n163) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n162) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n161) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n160) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n159) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n157) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n147) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n156) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n155) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n154) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n153) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n152) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n151) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n150) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n149) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n148) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n146) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n136) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n145) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n144) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n143) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n142) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n141) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n140) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n139) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n138) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n199) );
  INV_X1 U2 ( .A(c[10]), .ZN(n2) );
  INV_X1 U3 ( .A(a[10]), .ZN(n1) );
  INV_X1 U4 ( .A(a[7]), .ZN(n3) );
  XNOR2_X1 U5 ( .A(n1), .B(b[10]), .ZN(n137) );
  XNOR2_X1 U6 ( .A(n2), .B(n137), .ZN(result[10]) );
  XNOR2_X1 U7 ( .A(n3), .B(b[7]), .ZN(n197) );
  INV_X1 U8 ( .A(n24), .ZN(carry[28]) );
  AOI22_X1 U9 ( .A1(b[27]), .A2(a[27]), .B1(n155), .B2(c[27]), .ZN(n24) );
  INV_X1 U10 ( .A(n25), .ZN(carry[29]) );
  AOI22_X1 U11 ( .A1(b[28]), .A2(a[28]), .B1(n156), .B2(c[28]), .ZN(n25) );
  INV_X1 U12 ( .A(n27), .ZN(carry[30]) );
  AOI22_X1 U13 ( .A1(b[29]), .A2(a[29]), .B1(n157), .B2(c[29]), .ZN(n27) );
  INV_X1 U14 ( .A(n28), .ZN(carry[31]) );
  AOI22_X1 U15 ( .A1(b[30]), .A2(a[30]), .B1(n159), .B2(c[30]), .ZN(n28) );
  INV_X1 U16 ( .A(c[7]), .ZN(n4) );
  XOR2_X1 U17 ( .A(c[8]), .B(n198), .Z(result[8]) );
  INV_X1 U18 ( .A(n18), .ZN(carry[22]) );
  AOI22_X1 U19 ( .A1(b[21]), .A2(a[21]), .B1(n149), .B2(c[21]), .ZN(n18) );
  INV_X1 U20 ( .A(n16), .ZN(carry[20]) );
  AOI22_X1 U21 ( .A1(b[19]), .A2(a[19]), .B1(n146), .B2(c[19]), .ZN(n16) );
  INV_X1 U22 ( .A(n13), .ZN(carry[18]) );
  AOI22_X1 U23 ( .A1(b[17]), .A2(a[17]), .B1(n144), .B2(c[17]), .ZN(n13) );
  INV_X1 U24 ( .A(n17), .ZN(carry[21]) );
  AOI22_X1 U25 ( .A1(b[20]), .A2(a[20]), .B1(n148), .B2(c[20]), .ZN(n17) );
  INV_X1 U26 ( .A(n14), .ZN(carry[19]) );
  AOI22_X1 U27 ( .A1(b[18]), .A2(a[18]), .B1(n145), .B2(c[18]), .ZN(n14) );
  INV_X1 U28 ( .A(n11), .ZN(carry[16]) );
  AOI22_X1 U29 ( .A1(b[15]), .A2(a[15]), .B1(n142), .B2(c[15]), .ZN(n11) );
  INV_X1 U30 ( .A(n12), .ZN(carry[17]) );
  AOI22_X1 U31 ( .A1(b[16]), .A2(a[16]), .B1(n143), .B2(c[16]), .ZN(n12) );
  INV_X1 U32 ( .A(n19), .ZN(carry[23]) );
  AOI22_X1 U33 ( .A1(b[22]), .A2(a[22]), .B1(n150), .B2(c[22]), .ZN(n19) );
  INV_X1 U34 ( .A(n20), .ZN(carry[24]) );
  AOI22_X1 U35 ( .A1(b[23]), .A2(a[23]), .B1(n151), .B2(c[23]), .ZN(n20) );
  INV_X1 U36 ( .A(n21), .ZN(carry[25]) );
  AOI22_X1 U37 ( .A1(b[24]), .A2(a[24]), .B1(n152), .B2(c[24]), .ZN(n21) );
  INV_X1 U38 ( .A(n22), .ZN(carry[26]) );
  AOI22_X1 U39 ( .A1(b[25]), .A2(a[25]), .B1(n153), .B2(c[25]), .ZN(n22) );
  INV_X1 U40 ( .A(n23), .ZN(carry[27]) );
  AOI22_X1 U41 ( .A1(b[26]), .A2(a[26]), .B1(n154), .B2(c[26]), .ZN(n23) );
  INV_X1 U42 ( .A(n9), .ZN(carry[14]) );
  AOI22_X1 U43 ( .A1(b[13]), .A2(a[13]), .B1(n140), .B2(c[13]), .ZN(n9) );
  INV_X1 U44 ( .A(n10), .ZN(carry[15]) );
  AOI22_X1 U45 ( .A1(b[14]), .A2(a[14]), .B1(n141), .B2(c[14]), .ZN(n10) );
  INV_X1 U46 ( .A(n29), .ZN(carry[32]) );
  AOI22_X1 U47 ( .A1(b[31]), .A2(a[31]), .B1(n160), .B2(c[31]), .ZN(n29) );
  INV_X1 U48 ( .A(n30), .ZN(carry[33]) );
  AOI22_X1 U49 ( .A1(b[32]), .A2(a[32]), .B1(n161), .B2(c[32]), .ZN(n30) );
  INV_X1 U50 ( .A(n31), .ZN(carry[34]) );
  AOI22_X1 U51 ( .A1(b[33]), .A2(a[33]), .B1(n162), .B2(c[33]), .ZN(n31) );
  INV_X1 U52 ( .A(n32), .ZN(carry[35]) );
  AOI22_X1 U53 ( .A1(b[34]), .A2(a[34]), .B1(n163), .B2(c[34]), .ZN(n32) );
  INV_X1 U54 ( .A(n33), .ZN(carry[36]) );
  AOI22_X1 U55 ( .A1(b[35]), .A2(a[35]), .B1(n164), .B2(c[35]), .ZN(n33) );
  INV_X1 U56 ( .A(n34), .ZN(carry[37]) );
  AOI22_X1 U57 ( .A1(b[36]), .A2(a[36]), .B1(n165), .B2(c[36]), .ZN(n34) );
  INV_X1 U58 ( .A(n35), .ZN(carry[38]) );
  AOI22_X1 U59 ( .A1(b[37]), .A2(a[37]), .B1(n166), .B2(c[37]), .ZN(n35) );
  INV_X1 U60 ( .A(n36), .ZN(carry[39]) );
  AOI22_X1 U61 ( .A1(b[38]), .A2(a[38]), .B1(n167), .B2(c[38]), .ZN(n36) );
  INV_X1 U62 ( .A(n38), .ZN(carry[40]) );
  AOI22_X1 U63 ( .A1(b[39]), .A2(a[39]), .B1(n168), .B2(c[39]), .ZN(n38) );
  INV_X1 U64 ( .A(n39), .ZN(carry[41]) );
  AOI22_X1 U65 ( .A1(b[40]), .A2(a[40]), .B1(n170), .B2(c[40]), .ZN(n39) );
  INV_X1 U66 ( .A(n40), .ZN(carry[42]) );
  AOI22_X1 U67 ( .A1(b[41]), .A2(a[41]), .B1(n171), .B2(c[41]), .ZN(n40) );
  INV_X1 U68 ( .A(n41), .ZN(carry[43]) );
  AOI22_X1 U69 ( .A1(b[42]), .A2(a[42]), .B1(n172), .B2(c[42]), .ZN(n41) );
  INV_X1 U70 ( .A(n43), .ZN(carry[45]) );
  AOI22_X1 U71 ( .A1(b[44]), .A2(a[44]), .B1(n174), .B2(c[44]), .ZN(n43) );
  INV_X1 U72 ( .A(n45), .ZN(carry[47]) );
  AOI22_X1 U73 ( .A1(b[46]), .A2(a[46]), .B1(n176), .B2(c[46]), .ZN(n45) );
  INV_X1 U74 ( .A(n46), .ZN(carry[48]) );
  AOI22_X1 U75 ( .A1(b[47]), .A2(a[47]), .B1(n177), .B2(c[47]), .ZN(n46) );
  INV_X1 U76 ( .A(n49), .ZN(carry[50]) );
  AOI22_X1 U77 ( .A1(b[49]), .A2(a[49]), .B1(n179), .B2(c[49]), .ZN(n49) );
  INV_X1 U78 ( .A(n42), .ZN(carry[44]) );
  AOI22_X1 U79 ( .A1(b[43]), .A2(a[43]), .B1(n173), .B2(c[43]), .ZN(n42) );
  INV_X1 U80 ( .A(n44), .ZN(carry[46]) );
  AOI22_X1 U81 ( .A1(b[45]), .A2(a[45]), .B1(n175), .B2(c[45]), .ZN(n44) );
  INV_X1 U82 ( .A(n47), .ZN(carry[49]) );
  AOI22_X1 U83 ( .A1(b[48]), .A2(a[48]), .B1(n178), .B2(c[48]), .ZN(n47) );
  INV_X1 U84 ( .A(n50), .ZN(carry[51]) );
  AOI22_X1 U85 ( .A1(b[50]), .A2(a[50]), .B1(n181), .B2(c[50]), .ZN(n50) );
  INV_X1 U86 ( .A(n51), .ZN(carry[52]) );
  AOI22_X1 U87 ( .A1(b[51]), .A2(a[51]), .B1(n182), .B2(c[51]), .ZN(n51) );
  INV_X1 U88 ( .A(n52), .ZN(carry[53]) );
  AOI22_X1 U89 ( .A1(b[52]), .A2(a[52]), .B1(n183), .B2(c[52]), .ZN(n52) );
  INV_X1 U90 ( .A(n53), .ZN(carry[54]) );
  AOI22_X1 U91 ( .A1(b[53]), .A2(a[53]), .B1(n184), .B2(c[53]), .ZN(n53) );
  INV_X1 U92 ( .A(n54), .ZN(carry[55]) );
  AOI22_X1 U93 ( .A1(b[54]), .A2(a[54]), .B1(n185), .B2(c[54]), .ZN(n54) );
  INV_X1 U94 ( .A(n55), .ZN(carry[56]) );
  AOI22_X1 U95 ( .A1(b[55]), .A2(a[55]), .B1(n186), .B2(c[55]), .ZN(n55) );
  INV_X1 U96 ( .A(n56), .ZN(carry[57]) );
  AOI22_X1 U97 ( .A1(b[56]), .A2(a[56]), .B1(n187), .B2(c[56]), .ZN(n56) );
  INV_X1 U98 ( .A(n57), .ZN(carry[58]) );
  AOI22_X1 U99 ( .A1(b[57]), .A2(a[57]), .B1(n188), .B2(c[57]), .ZN(n57) );
  INV_X1 U100 ( .A(n58), .ZN(carry[59]) );
  AOI22_X1 U101 ( .A1(b[58]), .A2(a[58]), .B1(n189), .B2(c[58]), .ZN(n58) );
  INV_X1 U102 ( .A(n60), .ZN(carry[60]) );
  AOI22_X1 U103 ( .A1(b[59]), .A2(a[59]), .B1(n190), .B2(c[59]), .ZN(n60) );
  INV_X1 U104 ( .A(n61), .ZN(carry[61]) );
  AOI22_X1 U105 ( .A1(b[60]), .A2(a[60]), .B1(n192), .B2(c[60]), .ZN(n61) );
  INV_X1 U106 ( .A(n62), .ZN(carry[62]) );
  AOI22_X1 U107 ( .A1(b[61]), .A2(a[61]), .B1(n193), .B2(c[61]), .ZN(n62) );
  INV_X1 U108 ( .A(n134), .ZN(carry[8]) );
  INV_X1 U109 ( .A(n135), .ZN(carry[9]) );
  INV_X1 U110 ( .A(n5), .ZN(carry[10]) );
  AOI22_X1 U111 ( .A1(b[9]), .A2(a[9]), .B1(n199), .B2(c[9]), .ZN(n5) );
  INV_X1 U112 ( .A(n6), .ZN(carry[11]) );
  AOI22_X1 U113 ( .A1(b[10]), .A2(a[10]), .B1(n137), .B2(c[10]), .ZN(n6) );
  INV_X1 U114 ( .A(n7), .ZN(carry[12]) );
  AOI22_X1 U115 ( .A1(b[11]), .A2(a[11]), .B1(n138), .B2(c[11]), .ZN(n7) );
  INV_X1 U116 ( .A(n8), .ZN(carry[13]) );
  AOI22_X1 U117 ( .A1(b[12]), .A2(a[12]), .B1(n139), .B2(c[12]), .ZN(n8) );
  INV_X1 U118 ( .A(n132), .ZN(carry[6]) );
  AOI22_X1 U119 ( .A1(b[5]), .A2(a[5]), .B1(n191), .B2(c[5]), .ZN(n132) );
  INV_X1 U120 ( .A(n133), .ZN(carry[7]) );
  AOI22_X1 U121 ( .A1(b[6]), .A2(a[6]), .B1(n196), .B2(c[6]), .ZN(n133) );
  INV_X1 U122 ( .A(n59), .ZN(carry[5]) );
  AOI22_X1 U123 ( .A1(b[4]), .A2(a[4]), .B1(n180), .B2(c[4]), .ZN(n59) );
  INV_X1 U124 ( .A(n48), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n169), .B2(c[3]), .ZN(n48) );
  INV_X1 U126 ( .A(n63), .ZN(carry[63]) );
  AOI22_X1 U127 ( .A1(b[62]), .A2(a[62]), .B1(n194), .B2(c[62]), .ZN(n63) );
  INV_X1 U129 ( .A(n37), .ZN(carry[3]) );
  AOI22_X1 U130 ( .A1(b[2]), .A2(a[2]), .B1(n158), .B2(c[2]), .ZN(n37) );
  INV_X1 U191 ( .A(n26), .ZN(carry[2]) );
  AOI22_X1 U194 ( .A1(b[1]), .A2(a[1]), .B1(n147), .B2(c[1]), .ZN(n26) );
  INV_X1 U254 ( .A(n15), .ZN(carry[1]) );
  AOI22_X1 U256 ( .A1(b[0]), .A2(a[0]), .B1(n136), .B2(c[0]), .ZN(n15) );
  XNOR2_X1 U257 ( .A(n197), .B(n4), .ZN(result[7]) );
  AOI22_X1 U258 ( .A1(b[7]), .A2(a[7]), .B1(n197), .B2(c[7]), .ZN(n134) );
  AOI22_X1 U259 ( .A1(b[8]), .A2(a[8]), .B1(n198), .B2(c[8]), .ZN(n135) );
endmodule


module BWAdder_8 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(n213), .B(c[9]), .Z(result[9]) );
  XOR2_X1 U129 ( .A(n212), .B(c[8]), .Z(result[8]) );
  XOR2_X1 U130 ( .A(n211), .B(c[7]), .Z(result[7]) );
  XOR2_X1 U131 ( .A(n210), .B(c[6]), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n209), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n209) );
  XOR2_X1 U134 ( .A(c[62]), .B(n208), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n207), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n206), .Z(result[60]) );
  XOR2_X1 U137 ( .A(n205), .B(c[5]), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n204), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n203), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n202), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n201), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n200), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n199), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n198), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n197), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n196), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n195), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n1), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n193), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n192), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n191), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n190), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n189), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n188), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n187), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n186), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n185), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n184), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n183), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n182), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n181), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n180), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n179), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n178), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n177), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n176), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n175), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n174), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n173), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n172), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n171), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n170), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n169), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n168), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n167), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n166), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n165), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n164), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n163), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n162), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n161), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n160), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n159), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n158), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n157), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n156), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n155), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n154), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n153), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n152), .Z(result[11]) );
  XOR2_X1 U191 ( .A(n151), .B(c[10]), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n150), .Z(result[0]) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n208) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n207) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n206) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n204) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n194) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n203) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n202) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n201) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n200) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n199) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n198) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n197) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n196) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n195) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n193) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n183) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n192) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n191) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n190) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n189) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n188) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n187) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n186) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n185) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n184) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n182) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n172) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n181) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n180) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n179) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n178) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n177) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n176) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n175) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n174) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n173) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n171) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n161) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n170) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n169) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n168) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n167) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n166) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n165) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n164) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n163) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n162) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n160) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n150) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n159) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n158) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n157) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n156) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n155) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n154) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n153) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n152) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n151) );
  INV_X1 U2 ( .A(b[5]), .ZN(n8) );
  CLKBUF_X1 U3 ( .A(n194), .Z(n1) );
  CLKBUF_X1 U4 ( .A(a[8]), .Z(n2) );
  CLKBUF_X1 U5 ( .A(a[7]), .Z(n3) );
  INV_X1 U6 ( .A(b[7]), .ZN(n4) );
  INV_X1 U7 ( .A(b[8]), .ZN(n7) );
  INV_X1 U8 ( .A(b[9]), .ZN(n5) );
  XNOR2_X1 U9 ( .A(a[7]), .B(n4), .ZN(n211) );
  XNOR2_X1 U10 ( .A(a[9]), .B(n5), .ZN(n213) );
  CLKBUF_X1 U11 ( .A(a[6]), .Z(n6) );
  XNOR2_X1 U12 ( .A(a[8]), .B(n7), .ZN(n212) );
  XNOR2_X1 U13 ( .A(a[5]), .B(n8), .ZN(n205) );
  CLKBUF_X1 U14 ( .A(a[5]), .Z(n9) );
  INV_X1 U15 ( .A(n13), .ZN(carry[11]) );
  INV_X1 U16 ( .A(n12), .ZN(carry[10]) );
  INV_X1 U17 ( .A(n55), .ZN(carry[4]) );
  AOI22_X1 U18 ( .A1(b[3]), .A2(a[3]), .B1(n183), .B2(c[3]), .ZN(n55) );
  INV_X1 U19 ( .A(b[6]), .ZN(n11) );
  INV_X1 U20 ( .A(n149), .ZN(carry[9]) );
  INV_X1 U21 ( .A(n25), .ZN(carry[22]) );
  AOI22_X1 U22 ( .A1(b[21]), .A2(a[21]), .B1(n163), .B2(c[21]), .ZN(n25) );
  INV_X1 U23 ( .A(n14), .ZN(carry[12]) );
  AOI22_X1 U24 ( .A1(b[11]), .A2(a[11]), .B1(n152), .B2(c[11]), .ZN(n14) );
  INV_X1 U25 ( .A(n15), .ZN(carry[13]) );
  AOI22_X1 U26 ( .A1(b[12]), .A2(a[12]), .B1(n153), .B2(c[12]), .ZN(n15) );
  INV_X1 U27 ( .A(n24), .ZN(carry[21]) );
  AOI22_X1 U28 ( .A1(b[20]), .A2(a[20]), .B1(n162), .B2(c[20]), .ZN(n24) );
  INV_X1 U29 ( .A(n23), .ZN(carry[20]) );
  AOI22_X1 U30 ( .A1(b[19]), .A2(a[19]), .B1(n160), .B2(c[19]), .ZN(n23) );
  INV_X1 U31 ( .A(n16), .ZN(carry[14]) );
  AOI22_X1 U32 ( .A1(b[13]), .A2(a[13]), .B1(n154), .B2(c[13]), .ZN(n16) );
  INV_X1 U33 ( .A(n17), .ZN(carry[15]) );
  AOI22_X1 U34 ( .A1(b[14]), .A2(a[14]), .B1(n155), .B2(c[14]), .ZN(n17) );
  INV_X1 U35 ( .A(n20), .ZN(carry[18]) );
  AOI22_X1 U36 ( .A1(b[17]), .A2(a[17]), .B1(n158), .B2(c[17]), .ZN(n20) );
  INV_X1 U37 ( .A(n21), .ZN(carry[19]) );
  AOI22_X1 U38 ( .A1(b[18]), .A2(a[18]), .B1(n159), .B2(c[18]), .ZN(n21) );
  INV_X1 U39 ( .A(n18), .ZN(carry[16]) );
  AOI22_X1 U40 ( .A1(b[15]), .A2(a[15]), .B1(n156), .B2(c[15]), .ZN(n18) );
  INV_X1 U41 ( .A(n19), .ZN(carry[17]) );
  AOI22_X1 U42 ( .A1(b[16]), .A2(a[16]), .B1(n157), .B2(c[16]), .ZN(n19) );
  INV_X1 U43 ( .A(n26), .ZN(carry[23]) );
  AOI22_X1 U44 ( .A1(b[22]), .A2(a[22]), .B1(n164), .B2(c[22]), .ZN(n26) );
  INV_X1 U45 ( .A(n27), .ZN(carry[24]) );
  AOI22_X1 U46 ( .A1(b[23]), .A2(a[23]), .B1(n165), .B2(c[23]), .ZN(n27) );
  INV_X1 U47 ( .A(n28), .ZN(carry[25]) );
  AOI22_X1 U48 ( .A1(b[24]), .A2(a[24]), .B1(n166), .B2(c[24]), .ZN(n28) );
  INV_X1 U49 ( .A(n29), .ZN(carry[26]) );
  AOI22_X1 U50 ( .A1(b[25]), .A2(a[25]), .B1(n167), .B2(c[25]), .ZN(n29) );
  INV_X1 U51 ( .A(n30), .ZN(carry[27]) );
  AOI22_X1 U52 ( .A1(b[26]), .A2(a[26]), .B1(n168), .B2(c[26]), .ZN(n30) );
  INV_X1 U53 ( .A(n31), .ZN(carry[28]) );
  AOI22_X1 U54 ( .A1(b[27]), .A2(a[27]), .B1(n169), .B2(c[27]), .ZN(n31) );
  INV_X1 U55 ( .A(n32), .ZN(carry[29]) );
  AOI22_X1 U56 ( .A1(b[28]), .A2(a[28]), .B1(n170), .B2(c[28]), .ZN(n32) );
  INV_X1 U57 ( .A(n34), .ZN(carry[30]) );
  AOI22_X1 U58 ( .A1(b[29]), .A2(a[29]), .B1(n171), .B2(c[29]), .ZN(n34) );
  INV_X1 U59 ( .A(n35), .ZN(carry[31]) );
  AOI22_X1 U60 ( .A1(b[30]), .A2(a[30]), .B1(n173), .B2(c[30]), .ZN(n35) );
  INV_X1 U61 ( .A(n141), .ZN(carry[5]) );
  INV_X1 U62 ( .A(n36), .ZN(carry[32]) );
  AOI22_X1 U63 ( .A1(b[31]), .A2(a[31]), .B1(n174), .B2(c[31]), .ZN(n36) );
  INV_X1 U64 ( .A(n37), .ZN(carry[33]) );
  AOI22_X1 U65 ( .A1(b[32]), .A2(a[32]), .B1(n175), .B2(c[32]), .ZN(n37) );
  INV_X1 U66 ( .A(n38), .ZN(carry[34]) );
  AOI22_X1 U67 ( .A1(b[33]), .A2(a[33]), .B1(n176), .B2(c[33]), .ZN(n38) );
  INV_X1 U68 ( .A(n39), .ZN(carry[35]) );
  AOI22_X1 U69 ( .A1(b[34]), .A2(a[34]), .B1(n177), .B2(c[34]), .ZN(n39) );
  INV_X1 U70 ( .A(n40), .ZN(carry[36]) );
  AOI22_X1 U71 ( .A1(b[35]), .A2(a[35]), .B1(n178), .B2(c[35]), .ZN(n40) );
  INV_X1 U72 ( .A(n41), .ZN(carry[37]) );
  AOI22_X1 U73 ( .A1(b[36]), .A2(a[36]), .B1(n179), .B2(c[36]), .ZN(n41) );
  INV_X1 U74 ( .A(n42), .ZN(carry[38]) );
  AOI22_X1 U75 ( .A1(b[37]), .A2(a[37]), .B1(n180), .B2(c[37]), .ZN(n42) );
  INV_X1 U76 ( .A(n43), .ZN(carry[39]) );
  AOI22_X1 U77 ( .A1(b[38]), .A2(a[38]), .B1(n181), .B2(c[38]), .ZN(n43) );
  INV_X1 U78 ( .A(n45), .ZN(carry[40]) );
  AOI22_X1 U79 ( .A1(b[39]), .A2(a[39]), .B1(n182), .B2(c[39]), .ZN(n45) );
  INV_X1 U80 ( .A(n46), .ZN(carry[41]) );
  AOI22_X1 U81 ( .A1(b[40]), .A2(a[40]), .B1(n184), .B2(c[40]), .ZN(n46) );
  INV_X1 U82 ( .A(n47), .ZN(carry[42]) );
  AOI22_X1 U83 ( .A1(b[41]), .A2(a[41]), .B1(n185), .B2(c[41]), .ZN(n47) );
  INV_X1 U84 ( .A(n48), .ZN(carry[43]) );
  AOI22_X1 U85 ( .A1(b[42]), .A2(a[42]), .B1(n186), .B2(c[42]), .ZN(n48) );
  INV_X1 U86 ( .A(n49), .ZN(carry[44]) );
  AOI22_X1 U87 ( .A1(b[43]), .A2(a[43]), .B1(n187), .B2(c[43]), .ZN(n49) );
  INV_X1 U88 ( .A(n50), .ZN(carry[45]) );
  AOI22_X1 U89 ( .A1(b[44]), .A2(a[44]), .B1(n188), .B2(c[44]), .ZN(n50) );
  INV_X1 U90 ( .A(n51), .ZN(carry[46]) );
  AOI22_X1 U91 ( .A1(b[45]), .A2(a[45]), .B1(n189), .B2(c[45]), .ZN(n51) );
  INV_X1 U92 ( .A(n52), .ZN(carry[47]) );
  AOI22_X1 U93 ( .A1(b[46]), .A2(a[46]), .B1(n190), .B2(c[46]), .ZN(n52) );
  INV_X1 U94 ( .A(n53), .ZN(carry[48]) );
  AOI22_X1 U95 ( .A1(b[47]), .A2(a[47]), .B1(n191), .B2(c[47]), .ZN(n53) );
  INV_X1 U96 ( .A(n54), .ZN(carry[49]) );
  AOI22_X1 U97 ( .A1(b[48]), .A2(a[48]), .B1(n192), .B2(c[48]), .ZN(n54) );
  INV_X1 U98 ( .A(n56), .ZN(carry[50]) );
  AOI22_X1 U99 ( .A1(b[49]), .A2(a[49]), .B1(n193), .B2(c[49]), .ZN(n56) );
  INV_X1 U100 ( .A(n57), .ZN(carry[51]) );
  AOI22_X1 U101 ( .A1(b[50]), .A2(a[50]), .B1(n195), .B2(c[50]), .ZN(n57) );
  INV_X1 U102 ( .A(n58), .ZN(carry[52]) );
  AOI22_X1 U103 ( .A1(b[51]), .A2(a[51]), .B1(n196), .B2(c[51]), .ZN(n58) );
  INV_X1 U104 ( .A(n59), .ZN(carry[53]) );
  AOI22_X1 U105 ( .A1(b[52]), .A2(a[52]), .B1(n197), .B2(c[52]), .ZN(n59) );
  INV_X1 U106 ( .A(n60), .ZN(carry[54]) );
  AOI22_X1 U107 ( .A1(b[53]), .A2(a[53]), .B1(n198), .B2(c[53]), .ZN(n60) );
  INV_X1 U108 ( .A(n61), .ZN(carry[55]) );
  AOI22_X1 U109 ( .A1(b[54]), .A2(a[54]), .B1(n199), .B2(c[54]), .ZN(n61) );
  INV_X1 U110 ( .A(n62), .ZN(carry[56]) );
  AOI22_X1 U111 ( .A1(b[55]), .A2(a[55]), .B1(n200), .B2(c[55]), .ZN(n62) );
  AOI22_X1 U112 ( .A1(b[62]), .A2(a[62]), .B1(n208), .B2(c[62]), .ZN(n145) );
  INV_X1 U113 ( .A(n63), .ZN(carry[57]) );
  AOI22_X1 U114 ( .A1(b[56]), .A2(a[56]), .B1(n201), .B2(c[56]), .ZN(n63) );
  INV_X1 U115 ( .A(n139), .ZN(carry[58]) );
  AOI22_X1 U116 ( .A1(b[57]), .A2(a[57]), .B1(n202), .B2(c[57]), .ZN(n139) );
  INV_X1 U117 ( .A(n140), .ZN(carry[59]) );
  AOI22_X1 U118 ( .A1(b[58]), .A2(a[58]), .B1(n203), .B2(c[58]), .ZN(n140) );
  INV_X1 U119 ( .A(n142), .ZN(carry[60]) );
  AOI22_X1 U120 ( .A1(b[59]), .A2(a[59]), .B1(n204), .B2(c[59]), .ZN(n142) );
  INV_X1 U121 ( .A(n143), .ZN(carry[61]) );
  AOI22_X1 U122 ( .A1(b[60]), .A2(a[60]), .B1(n206), .B2(c[60]), .ZN(n143) );
  INV_X1 U123 ( .A(n144), .ZN(carry[62]) );
  AOI22_X1 U124 ( .A1(b[61]), .A2(a[61]), .B1(n207), .B2(c[61]), .ZN(n144) );
  INV_X1 U125 ( .A(n145), .ZN(carry[63]) );
  INV_X1 U126 ( .A(n44), .ZN(carry[3]) );
  AOI22_X1 U127 ( .A1(b[2]), .A2(a[2]), .B1(n172), .B2(c[2]), .ZN(n44) );
  INV_X1 U193 ( .A(n33), .ZN(carry[2]) );
  AOI22_X1 U194 ( .A1(b[1]), .A2(a[1]), .B1(n161), .B2(c[1]), .ZN(n33) );
  INV_X1 U195 ( .A(n22), .ZN(carry[1]) );
  AOI22_X1 U196 ( .A1(b[0]), .A2(a[0]), .B1(n150), .B2(c[0]), .ZN(n22) );
  INV_X1 U255 ( .A(n147), .ZN(carry[7]) );
  CLKBUF_X1 U256 ( .A(n212), .Z(n10) );
  AOI22_X1 U257 ( .A1(b[4]), .A2(a[4]), .B1(n194), .B2(c[4]), .ZN(n141) );
  AOI22_X1 U258 ( .A1(b[10]), .A2(a[10]), .B1(n151), .B2(c[10]), .ZN(n13) );
  XNOR2_X1 U259 ( .A(a[6]), .B(n11), .ZN(n210) );
  AOI22_X1 U260 ( .A1(b[9]), .A2(a[9]), .B1(n213), .B2(c[9]), .ZN(n12) );
  AOI22_X1 U261 ( .A1(b[5]), .A2(n9), .B1(n205), .B2(c[5]), .ZN(n146) );
  AOI22_X1 U262 ( .A1(b[7]), .A2(n3), .B1(n211), .B2(c[7]), .ZN(n148) );
  INV_X1 U263 ( .A(n148), .ZN(carry[8]) );
  AOI22_X1 U264 ( .A1(b[6]), .A2(n6), .B1(n210), .B2(c[6]), .ZN(n147) );
  INV_X1 U265 ( .A(n146), .ZN(carry[6]) );
  AOI22_X1 U266 ( .A1(b[8]), .A2(n2), .B1(n10), .B2(c[8]), .ZN(n149) );
endmodule


module BWAdder_9 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U3 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U4 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U5 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U6 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U7 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U8 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U9 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U10 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U11 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U12 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U13 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U14 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U15 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U16 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U17 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U18 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U19 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U20 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U21 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U22 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U23 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U24 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U25 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U26 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U27 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U28 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U29 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U30 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U31 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U32 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U33 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U34 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U35 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U36 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U37 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U38 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U39 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U40 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U41 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U42 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U43 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U44 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U45 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U46 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U47 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U48 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U49 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U50 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U51 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U52 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U53 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U54 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U55 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U56 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U57 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U58 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U59 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U60 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U61 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U62 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U63 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U64 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U65 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U66 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U67 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U68 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U69 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U70 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U71 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U72 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U73 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U74 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U75 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U76 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U77 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U78 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U79 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U80 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U81 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U82 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U83 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U84 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U85 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U86 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U87 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U88 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U89 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U90 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U91 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U92 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U93 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U94 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U95 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U96 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U97 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U98 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U99 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U100 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U101 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U102 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U103 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U104 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U105 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U106 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U107 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U108 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U109 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U110 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U111 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U112 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U113 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U114 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U115 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U116 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U117 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U118 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U119 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U120 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U121 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U122 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U123 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U124 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U125 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_10 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n197), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n196), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n195), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n194), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n193), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n193) );
  XOR2_X1 U134 ( .A(c[62]), .B(n192), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n191), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n190), .Z(result[60]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n188), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n187), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n186), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n185), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n184), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n183), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n182), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n181), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n180), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n179), .Z(result[50]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n177), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n176), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n175), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n174), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n173), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n172), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n171), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n170), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n169), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n168), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n167), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n166), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n165), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n164), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n163), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n162), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n161), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n160), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n159), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n158), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n157), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n156), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n155), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n154), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n153), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n152), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n151), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n150), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n149), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n148), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n147), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n146), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n145), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n144), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n143), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n142), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n141), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n140), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n139), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n138), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n137), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n136), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n135), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n134), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n196) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n195) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n194) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n189) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n192) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n191) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n190) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n188) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n187) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n186) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n185) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n184) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n183) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n182) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n181) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n180) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n179) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n177) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n167) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n176) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n175) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n174) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n173) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n172) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n171) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n170) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n169) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n168) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n166) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n156) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n165) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n164) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n163) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n162) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n161) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n160) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n159) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n158) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n157) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n155) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n145) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n154) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n153) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n152) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n151) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n150) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n149) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n148) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n147) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n146) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n144) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n134) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n143) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n142) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n141) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n140) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n139) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n138) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n137) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n136) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n135) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n197) );
  INV_X1 U2 ( .A(b[4]), .ZN(n2) );
  INV_X1 U3 ( .A(c[5]), .ZN(n3) );
  INV_X1 U4 ( .A(c[4]), .ZN(n1) );
  XNOR2_X1 U5 ( .A(n1), .B(n178), .ZN(result[4]) );
  XNOR2_X1 U6 ( .A(a[4]), .B(n2), .ZN(n178) );
  XNOR2_X1 U7 ( .A(n3), .B(n189), .ZN(result[5]) );
  INV_X1 U8 ( .A(n55), .ZN(carry[57]) );
  AOI22_X1 U9 ( .A1(b[56]), .A2(a[56]), .B1(n185), .B2(c[56]), .ZN(n55) );
  INV_X1 U10 ( .A(n61), .ZN(carry[62]) );
  AOI22_X1 U11 ( .A1(b[61]), .A2(a[61]), .B1(n191), .B2(c[61]), .ZN(n61) );
  INV_X1 U12 ( .A(n56), .ZN(carry[58]) );
  AOI22_X1 U13 ( .A1(b[57]), .A2(a[57]), .B1(n186), .B2(c[57]), .ZN(n56) );
  INV_X1 U14 ( .A(n57), .ZN(carry[59]) );
  AOI22_X1 U15 ( .A1(b[58]), .A2(a[58]), .B1(n187), .B2(c[58]), .ZN(n57) );
  INV_X1 U16 ( .A(n59), .ZN(carry[60]) );
  AOI22_X1 U17 ( .A1(b[59]), .A2(a[59]), .B1(n188), .B2(c[59]), .ZN(n59) );
  INV_X1 U18 ( .A(n60), .ZN(carry[61]) );
  AOI22_X1 U19 ( .A1(b[60]), .A2(a[60]), .B1(n190), .B2(c[60]), .ZN(n60) );
  INV_X1 U20 ( .A(n24), .ZN(carry[29]) );
  AOI22_X1 U21 ( .A1(b[28]), .A2(a[28]), .B1(n154), .B2(c[28]), .ZN(n24) );
  INV_X1 U22 ( .A(n26), .ZN(carry[30]) );
  AOI22_X1 U23 ( .A1(b[29]), .A2(a[29]), .B1(n155), .B2(c[29]), .ZN(n26) );
  INV_X1 U24 ( .A(n21), .ZN(carry[26]) );
  AOI22_X1 U25 ( .A1(b[25]), .A2(a[25]), .B1(n151), .B2(c[25]), .ZN(n21) );
  INV_X1 U26 ( .A(n22), .ZN(carry[27]) );
  AOI22_X1 U27 ( .A1(b[26]), .A2(a[26]), .B1(n152), .B2(c[26]), .ZN(n22) );
  INV_X1 U28 ( .A(n23), .ZN(carry[28]) );
  AOI22_X1 U29 ( .A1(b[27]), .A2(a[27]), .B1(n153), .B2(c[27]), .ZN(n23) );
  INV_X1 U30 ( .A(n19), .ZN(carry[24]) );
  AOI22_X1 U31 ( .A1(b[23]), .A2(a[23]), .B1(n149), .B2(c[23]), .ZN(n19) );
  INV_X1 U32 ( .A(n20), .ZN(carry[25]) );
  AOI22_X1 U33 ( .A1(b[24]), .A2(a[24]), .B1(n150), .B2(c[24]), .ZN(n20) );
  INV_X1 U34 ( .A(n17), .ZN(carry[22]) );
  AOI22_X1 U35 ( .A1(b[21]), .A2(a[21]), .B1(n147), .B2(c[21]), .ZN(n17) );
  INV_X1 U36 ( .A(n18), .ZN(carry[23]) );
  AOI22_X1 U37 ( .A1(b[22]), .A2(a[22]), .B1(n148), .B2(c[22]), .ZN(n18) );
  INV_X1 U38 ( .A(n27), .ZN(carry[31]) );
  AOI22_X1 U39 ( .A1(b[30]), .A2(a[30]), .B1(n157), .B2(c[30]), .ZN(n27) );
  INV_X1 U40 ( .A(n28), .ZN(carry[32]) );
  AOI22_X1 U41 ( .A1(b[31]), .A2(a[31]), .B1(n158), .B2(c[31]), .ZN(n28) );
  INV_X1 U42 ( .A(n29), .ZN(carry[33]) );
  AOI22_X1 U43 ( .A1(b[32]), .A2(a[32]), .B1(n159), .B2(c[32]), .ZN(n29) );
  INV_X1 U44 ( .A(n30), .ZN(carry[34]) );
  AOI22_X1 U45 ( .A1(b[33]), .A2(a[33]), .B1(n160), .B2(c[33]), .ZN(n30) );
  INV_X1 U46 ( .A(n31), .ZN(carry[35]) );
  AOI22_X1 U47 ( .A1(b[34]), .A2(a[34]), .B1(n161), .B2(c[34]), .ZN(n31) );
  INV_X1 U48 ( .A(n32), .ZN(carry[36]) );
  AOI22_X1 U49 ( .A1(b[35]), .A2(a[35]), .B1(n162), .B2(c[35]), .ZN(n32) );
  INV_X1 U50 ( .A(n33), .ZN(carry[37]) );
  AOI22_X1 U51 ( .A1(b[36]), .A2(a[36]), .B1(n163), .B2(c[36]), .ZN(n33) );
  INV_X1 U52 ( .A(n34), .ZN(carry[38]) );
  AOI22_X1 U53 ( .A1(b[37]), .A2(a[37]), .B1(n164), .B2(c[37]), .ZN(n34) );
  INV_X1 U54 ( .A(n35), .ZN(carry[39]) );
  AOI22_X1 U55 ( .A1(b[38]), .A2(a[38]), .B1(n165), .B2(c[38]), .ZN(n35) );
  INV_X1 U56 ( .A(n37), .ZN(carry[40]) );
  AOI22_X1 U57 ( .A1(b[39]), .A2(a[39]), .B1(n166), .B2(c[39]), .ZN(n37) );
  INV_X1 U58 ( .A(n38), .ZN(carry[41]) );
  AOI22_X1 U59 ( .A1(b[40]), .A2(a[40]), .B1(n168), .B2(c[40]), .ZN(n38) );
  INV_X1 U60 ( .A(n39), .ZN(carry[42]) );
  AOI22_X1 U61 ( .A1(b[41]), .A2(a[41]), .B1(n169), .B2(c[41]), .ZN(n39) );
  INV_X1 U62 ( .A(n40), .ZN(carry[43]) );
  AOI22_X1 U63 ( .A1(b[42]), .A2(a[42]), .B1(n170), .B2(c[42]), .ZN(n40) );
  INV_X1 U64 ( .A(n41), .ZN(carry[44]) );
  AOI22_X1 U65 ( .A1(b[43]), .A2(a[43]), .B1(n171), .B2(c[43]), .ZN(n41) );
  INV_X1 U66 ( .A(n42), .ZN(carry[45]) );
  AOI22_X1 U67 ( .A1(b[44]), .A2(a[44]), .B1(n172), .B2(c[44]), .ZN(n42) );
  INV_X1 U68 ( .A(n46), .ZN(carry[49]) );
  AOI22_X1 U69 ( .A1(b[48]), .A2(a[48]), .B1(n176), .B2(c[48]), .ZN(n46) );
  INV_X1 U70 ( .A(n49), .ZN(carry[51]) );
  AOI22_X1 U71 ( .A1(b[50]), .A2(a[50]), .B1(n179), .B2(c[50]), .ZN(n49) );
  INV_X1 U72 ( .A(n50), .ZN(carry[52]) );
  AOI22_X1 U73 ( .A1(b[51]), .A2(a[51]), .B1(n180), .B2(c[51]), .ZN(n50) );
  INV_X1 U74 ( .A(n52), .ZN(carry[54]) );
  AOI22_X1 U75 ( .A1(b[53]), .A2(a[53]), .B1(n182), .B2(c[53]), .ZN(n52) );
  INV_X1 U76 ( .A(n53), .ZN(carry[55]) );
  AOI22_X1 U77 ( .A1(b[54]), .A2(a[54]), .B1(n183), .B2(c[54]), .ZN(n53) );
  INV_X1 U78 ( .A(n43), .ZN(carry[46]) );
  AOI22_X1 U79 ( .A1(b[45]), .A2(a[45]), .B1(n173), .B2(c[45]), .ZN(n43) );
  INV_X1 U80 ( .A(n44), .ZN(carry[47]) );
  AOI22_X1 U81 ( .A1(b[46]), .A2(a[46]), .B1(n174), .B2(c[46]), .ZN(n44) );
  INV_X1 U82 ( .A(n45), .ZN(carry[48]) );
  AOI22_X1 U83 ( .A1(b[47]), .A2(a[47]), .B1(n175), .B2(c[47]), .ZN(n45) );
  INV_X1 U84 ( .A(n48), .ZN(carry[50]) );
  AOI22_X1 U85 ( .A1(b[49]), .A2(a[49]), .B1(n177), .B2(c[49]), .ZN(n48) );
  INV_X1 U86 ( .A(n51), .ZN(carry[53]) );
  AOI22_X1 U87 ( .A1(b[52]), .A2(a[52]), .B1(n181), .B2(c[52]), .ZN(n51) );
  INV_X1 U88 ( .A(n54), .ZN(carry[56]) );
  AOI22_X1 U89 ( .A1(b[55]), .A2(a[55]), .B1(n184), .B2(c[55]), .ZN(n54) );
  INV_X1 U90 ( .A(n58), .ZN(carry[5]) );
  INV_X1 U91 ( .A(n63), .ZN(carry[6]) );
  INV_X1 U92 ( .A(n47), .ZN(carry[4]) );
  AOI22_X1 U93 ( .A1(b[3]), .A2(a[3]), .B1(n167), .B2(c[3]), .ZN(n47) );
  INV_X1 U94 ( .A(n131), .ZN(carry[7]) );
  AOI22_X1 U95 ( .A1(b[6]), .A2(a[6]), .B1(n194), .B2(c[6]), .ZN(n131) );
  INV_X1 U96 ( .A(n132), .ZN(carry[8]) );
  AOI22_X1 U97 ( .A1(b[7]), .A2(a[7]), .B1(n195), .B2(c[7]), .ZN(n132) );
  INV_X1 U98 ( .A(n133), .ZN(carry[9]) );
  AOI22_X1 U99 ( .A1(b[8]), .A2(a[8]), .B1(n196), .B2(c[8]), .ZN(n133) );
  INV_X1 U100 ( .A(n4), .ZN(carry[10]) );
  AOI22_X1 U101 ( .A1(b[9]), .A2(a[9]), .B1(n197), .B2(c[9]), .ZN(n4) );
  INV_X1 U102 ( .A(n5), .ZN(carry[11]) );
  AOI22_X1 U103 ( .A1(b[10]), .A2(a[10]), .B1(n135), .B2(c[10]), .ZN(n5) );
  INV_X1 U104 ( .A(n6), .ZN(carry[12]) );
  AOI22_X1 U105 ( .A1(b[11]), .A2(a[11]), .B1(n136), .B2(c[11]), .ZN(n6) );
  INV_X1 U106 ( .A(n7), .ZN(carry[13]) );
  AOI22_X1 U107 ( .A1(b[12]), .A2(a[12]), .B1(n137), .B2(c[12]), .ZN(n7) );
  INV_X1 U108 ( .A(n8), .ZN(carry[14]) );
  AOI22_X1 U109 ( .A1(b[13]), .A2(a[13]), .B1(n138), .B2(c[13]), .ZN(n8) );
  INV_X1 U110 ( .A(n9), .ZN(carry[15]) );
  AOI22_X1 U111 ( .A1(b[14]), .A2(a[14]), .B1(n139), .B2(c[14]), .ZN(n9) );
  INV_X1 U112 ( .A(n10), .ZN(carry[16]) );
  AOI22_X1 U113 ( .A1(b[15]), .A2(a[15]), .B1(n140), .B2(c[15]), .ZN(n10) );
  INV_X1 U114 ( .A(n11), .ZN(carry[17]) );
  AOI22_X1 U115 ( .A1(b[16]), .A2(a[16]), .B1(n141), .B2(c[16]), .ZN(n11) );
  INV_X1 U116 ( .A(n12), .ZN(carry[18]) );
  AOI22_X1 U117 ( .A1(b[17]), .A2(a[17]), .B1(n142), .B2(c[17]), .ZN(n12) );
  INV_X1 U118 ( .A(n13), .ZN(carry[19]) );
  AOI22_X1 U119 ( .A1(b[18]), .A2(a[18]), .B1(n143), .B2(c[18]), .ZN(n13) );
  INV_X1 U120 ( .A(n15), .ZN(carry[20]) );
  AOI22_X1 U121 ( .A1(b[19]), .A2(a[19]), .B1(n144), .B2(c[19]), .ZN(n15) );
  INV_X1 U122 ( .A(n16), .ZN(carry[21]) );
  AOI22_X1 U123 ( .A1(b[20]), .A2(a[20]), .B1(n146), .B2(c[20]), .ZN(n16) );
  INV_X1 U124 ( .A(n36), .ZN(carry[3]) );
  AOI22_X1 U125 ( .A1(b[2]), .A2(a[2]), .B1(n156), .B2(c[2]), .ZN(n36) );
  INV_X1 U126 ( .A(n62), .ZN(carry[63]) );
  AOI22_X1 U127 ( .A1(b[62]), .A2(a[62]), .B1(n192), .B2(c[62]), .ZN(n62) );
  INV_X1 U137 ( .A(n25), .ZN(carry[2]) );
  AOI22_X1 U148 ( .A1(b[1]), .A2(a[1]), .B1(n145), .B2(c[1]), .ZN(n25) );
  INV_X1 U201 ( .A(n14), .ZN(carry[1]) );
  AOI22_X1 U256 ( .A1(b[0]), .A2(a[0]), .B1(n134), .B2(c[0]), .ZN(n14) );
  AOI22_X1 U257 ( .A1(b[4]), .A2(a[4]), .B1(n178), .B2(c[4]), .ZN(n58) );
  AOI22_X1 U258 ( .A1(b[5]), .A2(a[5]), .B1(n189), .B2(c[5]), .ZN(n63) );
endmodule


module BWAdder_11 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  XOR2_X1 U2 ( .A(c[5]), .B(n183), .Z(result[5]) );
  INV_X1 U3 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U4 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U5 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U6 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U7 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U8 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U9 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U10 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U11 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U12 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U13 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U14 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U15 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U16 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U17 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U18 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U19 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U20 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U21 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U22 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U23 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U24 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U25 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U26 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U27 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U28 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U29 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U30 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U31 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U32 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U33 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U34 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U35 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U36 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U37 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U38 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U39 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U40 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U41 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U42 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U43 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U44 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U45 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U46 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U47 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U48 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U49 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U50 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U51 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U52 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U53 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U54 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U55 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U56 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U57 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U58 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U59 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U60 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U61 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U62 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U63 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U64 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U65 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U66 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U67 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U68 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U69 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U70 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U71 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U72 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U73 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U74 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U75 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U76 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U77 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U78 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U79 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U80 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U81 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U82 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U83 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U84 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U85 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U86 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U87 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U88 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U89 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U90 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U91 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U92 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U93 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U94 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U95 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U96 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U97 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U98 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U99 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U100 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U101 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U102 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U103 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U104 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U105 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U106 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U107 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U108 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U109 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U110 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U111 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U112 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U113 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U114 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U115 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U116 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U117 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U118 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U119 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U120 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U121 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U122 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U123 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U124 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U125 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U126 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U127 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U137 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_12 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(n217), .B(c[9]), .Z(result[9]) );
  XOR2_X1 U129 ( .A(n216), .B(c[8]), .Z(result[8]) );
  XOR2_X1 U130 ( .A(n215), .B(c[7]), .Z(result[7]) );
  XOR2_X1 U131 ( .A(n214), .B(c[6]), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n213), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n213) );
  XOR2_X1 U134 ( .A(c[62]), .B(n212), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n211), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n210), .Z(result[60]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n208), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n207), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n206), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n205), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n204), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n203), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n202), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n201), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n200), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n199), .Z(result[50]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n197), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n196), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n195), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n194), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n193), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n192), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n191), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n190), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n189), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n188), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n187), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n186), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n185), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n184), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n183), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n182), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n181), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n180), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n179), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n178), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n177), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n176), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n175), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n174), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n173), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n172), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n171), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n170), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n169), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n168), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n167), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n166), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n165), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n164), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n163), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n162), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n161), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n160), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n159), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n158), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n157), .Z(result[12]) );
  XOR2_X1 U190 ( .A(n156), .B(c[11]), .Z(result[11]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n154), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n216) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n215) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n214) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n209) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n212) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n211) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n210) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n208) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n198) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n207) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n206) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n205) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n204) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n203) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n202) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n201) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n200) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n199) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n197) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n187) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n196) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n195) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n194) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n193) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n192) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n191) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n190) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n189) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n188) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n186) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n176) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n185) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n184) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n183) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n182) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n181) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n180) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n179) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n178) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n177) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n175) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n165) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n174) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n173) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n172) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n171) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n170) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n169) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n168) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n167) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n166) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n164) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n154) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n163) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n162) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n161) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n160) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n159) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n158) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n157) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n156) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n155) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n217) );
  CLKBUF_X1 U2 ( .A(a[10]), .Z(n1) );
  XOR2_X1 U3 ( .A(a[7]), .B(b[7]), .Z(n2) );
  XNOR2_X1 U4 ( .A(a[10]), .B(b[10]), .ZN(n3) );
  INV_X1 U5 ( .A(c[4]), .ZN(n10) );
  INV_X1 U6 ( .A(c[5]), .ZN(n11) );
  CLKBUF_X1 U7 ( .A(a[5]), .Z(n4) );
  CLKBUF_X1 U8 ( .A(a[9]), .Z(n5) );
  CLKBUF_X1 U9 ( .A(a[6]), .Z(n6) );
  NAND2_X1 U10 ( .A1(c[10]), .A2(n3), .ZN(n8) );
  NAND2_X1 U11 ( .A1(n7), .A2(n155), .ZN(n9) );
  NAND2_X1 U12 ( .A1(n8), .A2(n9), .ZN(result[10]) );
  INV_X1 U13 ( .A(c[10]), .ZN(n7) );
  XNOR2_X1 U14 ( .A(n10), .B(n198), .ZN(result[4]) );
  XNOR2_X1 U15 ( .A(n209), .B(n11), .ZN(result[5]) );
  INV_X1 U16 ( .A(n141), .ZN(carry[56]) );
  AOI22_X1 U17 ( .A1(b[55]), .A2(a[55]), .B1(n204), .B2(c[55]), .ZN(n141) );
  INV_X1 U18 ( .A(n142), .ZN(carry[57]) );
  AOI22_X1 U19 ( .A1(b[56]), .A2(a[56]), .B1(n205), .B2(c[56]), .ZN(n142) );
  INV_X1 U20 ( .A(n143), .ZN(carry[58]) );
  AOI22_X1 U21 ( .A1(b[57]), .A2(a[57]), .B1(n206), .B2(c[57]), .ZN(n143) );
  INV_X1 U22 ( .A(n144), .ZN(carry[59]) );
  AOI22_X1 U23 ( .A1(b[58]), .A2(a[58]), .B1(n207), .B2(c[58]), .ZN(n144) );
  INV_X1 U24 ( .A(n146), .ZN(carry[60]) );
  AOI22_X1 U25 ( .A1(b[59]), .A2(a[59]), .B1(n208), .B2(c[59]), .ZN(n146) );
  INV_X1 U26 ( .A(n147), .ZN(carry[61]) );
  AOI22_X1 U27 ( .A1(b[60]), .A2(a[60]), .B1(n210), .B2(c[60]), .ZN(n147) );
  INV_X1 U28 ( .A(n148), .ZN(carry[62]) );
  AOI22_X1 U29 ( .A1(b[61]), .A2(a[61]), .B1(n211), .B2(c[61]), .ZN(n148) );
  INV_X1 U30 ( .A(n149), .ZN(carry[63]) );
  AOI22_X1 U31 ( .A1(b[62]), .A2(a[62]), .B1(n212), .B2(c[62]), .ZN(n149) );
  INV_X1 U32 ( .A(n16), .ZN(carry[12]) );
  AOI22_X1 U33 ( .A1(b[11]), .A2(a[11]), .B1(n156), .B2(c[11]), .ZN(n16) );
  INV_X1 U34 ( .A(n17), .ZN(carry[13]) );
  AOI22_X1 U35 ( .A1(b[12]), .A2(a[12]), .B1(n157), .B2(c[12]), .ZN(n17) );
  INV_X1 U36 ( .A(n18), .ZN(carry[14]) );
  AOI22_X1 U37 ( .A1(b[13]), .A2(a[13]), .B1(n158), .B2(c[13]), .ZN(n18) );
  INV_X1 U38 ( .A(n19), .ZN(carry[15]) );
  AOI22_X1 U39 ( .A1(b[14]), .A2(a[14]), .B1(n159), .B2(c[14]), .ZN(n19) );
  INV_X1 U40 ( .A(n20), .ZN(carry[16]) );
  AOI22_X1 U41 ( .A1(b[15]), .A2(a[15]), .B1(n160), .B2(c[15]), .ZN(n20) );
  INV_X1 U42 ( .A(n36), .ZN(carry[30]) );
  AOI22_X1 U43 ( .A1(b[29]), .A2(a[29]), .B1(n175), .B2(c[29]), .ZN(n36) );
  INV_X1 U44 ( .A(n37), .ZN(carry[31]) );
  AOI22_X1 U45 ( .A1(b[30]), .A2(a[30]), .B1(n177), .B2(c[30]), .ZN(n37) );
  INV_X1 U46 ( .A(n15), .ZN(carry[11]) );
  AOI22_X1 U47 ( .A1(b[10]), .A2(n1), .B1(n155), .B2(c[10]), .ZN(n15) );
  INV_X1 U48 ( .A(n153), .ZN(carry[9]) );
  INV_X1 U49 ( .A(n14), .ZN(carry[10]) );
  INV_X1 U50 ( .A(n150), .ZN(carry[6]) );
  INV_X1 U51 ( .A(n145), .ZN(carry[5]) );
  INV_X1 U52 ( .A(n27), .ZN(carry[22]) );
  AOI22_X1 U53 ( .A1(b[21]), .A2(a[21]), .B1(n167), .B2(c[21]), .ZN(n27) );
  INV_X1 U54 ( .A(n26), .ZN(carry[21]) );
  AOI22_X1 U55 ( .A1(b[20]), .A2(a[20]), .B1(n166), .B2(c[20]), .ZN(n26) );
  INV_X1 U56 ( .A(n25), .ZN(carry[20]) );
  AOI22_X1 U57 ( .A1(b[19]), .A2(a[19]), .B1(n164), .B2(c[19]), .ZN(n25) );
  INV_X1 U58 ( .A(n22), .ZN(carry[18]) );
  AOI22_X1 U59 ( .A1(b[17]), .A2(a[17]), .B1(n162), .B2(c[17]), .ZN(n22) );
  INV_X1 U60 ( .A(n23), .ZN(carry[19]) );
  AOI22_X1 U61 ( .A1(b[18]), .A2(a[18]), .B1(n163), .B2(c[18]), .ZN(n23) );
  INV_X1 U62 ( .A(n21), .ZN(carry[17]) );
  AOI22_X1 U63 ( .A1(b[16]), .A2(a[16]), .B1(n161), .B2(c[16]), .ZN(n21) );
  INV_X1 U64 ( .A(n28), .ZN(carry[23]) );
  AOI22_X1 U65 ( .A1(b[22]), .A2(a[22]), .B1(n168), .B2(c[22]), .ZN(n28) );
  INV_X1 U66 ( .A(n29), .ZN(carry[24]) );
  AOI22_X1 U67 ( .A1(b[23]), .A2(a[23]), .B1(n169), .B2(c[23]), .ZN(n29) );
  INV_X1 U68 ( .A(n30), .ZN(carry[25]) );
  AOI22_X1 U69 ( .A1(b[24]), .A2(a[24]), .B1(n170), .B2(c[24]), .ZN(n30) );
  INV_X1 U70 ( .A(n31), .ZN(carry[26]) );
  AOI22_X1 U71 ( .A1(b[25]), .A2(a[25]), .B1(n171), .B2(c[25]), .ZN(n31) );
  INV_X1 U72 ( .A(n32), .ZN(carry[27]) );
  AOI22_X1 U73 ( .A1(b[26]), .A2(a[26]), .B1(n172), .B2(c[26]), .ZN(n32) );
  INV_X1 U74 ( .A(n33), .ZN(carry[28]) );
  AOI22_X1 U75 ( .A1(b[27]), .A2(a[27]), .B1(n173), .B2(c[27]), .ZN(n33) );
  INV_X1 U76 ( .A(n34), .ZN(carry[29]) );
  AOI22_X1 U77 ( .A1(b[28]), .A2(a[28]), .B1(n174), .B2(c[28]), .ZN(n34) );
  INV_X1 U78 ( .A(n152), .ZN(carry[8]) );
  INV_X1 U79 ( .A(n38), .ZN(carry[32]) );
  AOI22_X1 U80 ( .A1(b[31]), .A2(a[31]), .B1(n178), .B2(c[31]), .ZN(n38) );
  INV_X1 U81 ( .A(n39), .ZN(carry[33]) );
  AOI22_X1 U82 ( .A1(b[32]), .A2(a[32]), .B1(n179), .B2(c[32]), .ZN(n39) );
  INV_X1 U83 ( .A(n40), .ZN(carry[34]) );
  AOI22_X1 U84 ( .A1(b[33]), .A2(a[33]), .B1(n180), .B2(c[33]), .ZN(n40) );
  INV_X1 U85 ( .A(n41), .ZN(carry[35]) );
  AOI22_X1 U86 ( .A1(b[34]), .A2(a[34]), .B1(n181), .B2(c[34]), .ZN(n41) );
  INV_X1 U87 ( .A(n42), .ZN(carry[36]) );
  AOI22_X1 U88 ( .A1(b[35]), .A2(a[35]), .B1(n182), .B2(c[35]), .ZN(n42) );
  INV_X1 U89 ( .A(n43), .ZN(carry[37]) );
  AOI22_X1 U90 ( .A1(b[36]), .A2(a[36]), .B1(n183), .B2(c[36]), .ZN(n43) );
  INV_X1 U91 ( .A(n44), .ZN(carry[38]) );
  AOI22_X1 U92 ( .A1(b[37]), .A2(a[37]), .B1(n184), .B2(c[37]), .ZN(n44) );
  INV_X1 U93 ( .A(n45), .ZN(carry[39]) );
  AOI22_X1 U94 ( .A1(b[38]), .A2(a[38]), .B1(n185), .B2(c[38]), .ZN(n45) );
  INV_X1 U95 ( .A(n47), .ZN(carry[40]) );
  AOI22_X1 U96 ( .A1(b[39]), .A2(a[39]), .B1(n186), .B2(c[39]), .ZN(n47) );
  INV_X1 U97 ( .A(n48), .ZN(carry[41]) );
  AOI22_X1 U98 ( .A1(b[40]), .A2(a[40]), .B1(n188), .B2(c[40]), .ZN(n48) );
  INV_X1 U99 ( .A(n49), .ZN(carry[42]) );
  AOI22_X1 U100 ( .A1(b[41]), .A2(a[41]), .B1(n189), .B2(c[41]), .ZN(n49) );
  INV_X1 U101 ( .A(n50), .ZN(carry[43]) );
  AOI22_X1 U102 ( .A1(b[42]), .A2(a[42]), .B1(n190), .B2(c[42]), .ZN(n50) );
  INV_X1 U103 ( .A(n51), .ZN(carry[44]) );
  AOI22_X1 U104 ( .A1(b[43]), .A2(a[43]), .B1(n191), .B2(c[43]), .ZN(n51) );
  INV_X1 U105 ( .A(n55), .ZN(carry[48]) );
  AOI22_X1 U106 ( .A1(b[47]), .A2(a[47]), .B1(n195), .B2(c[47]), .ZN(n55) );
  INV_X1 U107 ( .A(n52), .ZN(carry[45]) );
  AOI22_X1 U108 ( .A1(b[44]), .A2(a[44]), .B1(n192), .B2(c[44]), .ZN(n52) );
  INV_X1 U109 ( .A(n53), .ZN(carry[46]) );
  AOI22_X1 U110 ( .A1(b[45]), .A2(a[45]), .B1(n193), .B2(c[45]), .ZN(n53) );
  INV_X1 U111 ( .A(n54), .ZN(carry[47]) );
  AOI22_X1 U112 ( .A1(b[46]), .A2(a[46]), .B1(n194), .B2(c[46]), .ZN(n54) );
  INV_X1 U113 ( .A(n56), .ZN(carry[49]) );
  AOI22_X1 U114 ( .A1(b[48]), .A2(a[48]), .B1(n196), .B2(c[48]), .ZN(n56) );
  INV_X1 U115 ( .A(n58), .ZN(carry[50]) );
  AOI22_X1 U116 ( .A1(b[49]), .A2(a[49]), .B1(n197), .B2(c[49]), .ZN(n58) );
  INV_X1 U117 ( .A(n59), .ZN(carry[51]) );
  AOI22_X1 U118 ( .A1(b[50]), .A2(a[50]), .B1(n199), .B2(c[50]), .ZN(n59) );
  INV_X1 U119 ( .A(n60), .ZN(carry[52]) );
  AOI22_X1 U120 ( .A1(b[51]), .A2(a[51]), .B1(n200), .B2(c[51]), .ZN(n60) );
  INV_X1 U121 ( .A(n61), .ZN(carry[53]) );
  AOI22_X1 U122 ( .A1(b[52]), .A2(a[52]), .B1(n201), .B2(c[52]), .ZN(n61) );
  INV_X1 U123 ( .A(n62), .ZN(carry[54]) );
  AOI22_X1 U124 ( .A1(b[53]), .A2(a[53]), .B1(n202), .B2(c[53]), .ZN(n62) );
  INV_X1 U125 ( .A(n63), .ZN(carry[55]) );
  AOI22_X1 U126 ( .A1(b[54]), .A2(a[54]), .B1(n203), .B2(c[54]), .ZN(n63) );
  INV_X1 U127 ( .A(n46), .ZN(carry[3]) );
  AOI22_X1 U137 ( .A1(b[2]), .A2(a[2]), .B1(n176), .B2(c[2]), .ZN(n46) );
  INV_X1 U148 ( .A(n57), .ZN(carry[4]) );
  AOI22_X1 U191 ( .A1(b[3]), .A2(a[3]), .B1(n187), .B2(c[3]), .ZN(n57) );
  INV_X1 U256 ( .A(n35), .ZN(carry[2]) );
  AOI22_X1 U257 ( .A1(b[1]), .A2(a[1]), .B1(n165), .B2(c[1]), .ZN(n35) );
  INV_X1 U258 ( .A(n24), .ZN(carry[1]) );
  AOI22_X1 U259 ( .A1(b[0]), .A2(a[0]), .B1(n154), .B2(c[0]), .ZN(n24) );
  INV_X1 U260 ( .A(n151), .ZN(carry[7]) );
  CLKBUF_X1 U261 ( .A(b[7]), .Z(n12) );
  CLKBUF_X1 U262 ( .A(a[8]), .Z(n13) );
  AOI22_X1 U263 ( .A1(b[9]), .A2(n5), .B1(n217), .B2(c[9]), .ZN(n14) );
  AOI22_X1 U264 ( .A1(b[4]), .A2(a[4]), .B1(n198), .B2(c[4]), .ZN(n145) );
  AOI22_X1 U265 ( .A1(b[5]), .A2(n4), .B1(n209), .B2(c[5]), .ZN(n150) );
  AOI22_X1 U266 ( .A1(b[6]), .A2(n6), .B1(n214), .B2(c[6]), .ZN(n151) );
  AOI22_X1 U267 ( .A1(n12), .A2(a[7]), .B1(n2), .B2(c[7]), .ZN(n152) );
  AOI22_X1 U268 ( .A1(b[8]), .A2(n13), .B1(n216), .B2(c[8]), .ZN(n153) );
endmodule


module BWAdder_13 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n59), .ZN(carry[63]) );
  INV_X1 U3 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U4 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U5 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U6 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U7 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U8 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U9 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U10 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U11 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U12 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U13 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U14 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U15 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U16 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U17 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U18 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U19 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U20 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U21 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U22 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U23 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U24 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U25 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U26 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U27 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U28 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U29 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U30 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U31 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U32 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U33 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U34 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U35 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U36 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U37 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U38 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U39 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U40 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U41 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U42 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U43 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U44 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  AOI22_X1 U45 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U46 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U47 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U48 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U49 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U50 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U51 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U52 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U53 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U54 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U55 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U56 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U57 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U58 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U59 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U60 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U61 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U62 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U63 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U64 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U65 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U66 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U67 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U68 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U69 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U70 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U71 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U72 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U73 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U74 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U75 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U76 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U77 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U78 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U79 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U80 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U81 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U82 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U83 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U84 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U85 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U86 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U87 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U88 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U89 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U90 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U91 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U92 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U93 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U94 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U95 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U96 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U97 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U98 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U99 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U100 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U101 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U102 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U103 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U104 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U105 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U106 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U107 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U108 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U109 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U110 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U111 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U112 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U113 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U114 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U115 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U116 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U117 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U118 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U119 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U120 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U121 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U122 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U123 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U124 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U125 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_14 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U3 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U4 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U5 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U6 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U7 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U8 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U9 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U10 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U11 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U12 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U13 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U14 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U15 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U16 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U17 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U18 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U19 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U20 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U21 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U22 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U23 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U24 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U25 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U26 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U27 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U28 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U29 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U30 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U31 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U32 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U33 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U34 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U35 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U36 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U37 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U38 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U39 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U40 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U41 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U42 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U43 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U44 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U45 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U46 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U47 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U48 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U49 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U50 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U51 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U52 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U53 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U54 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U55 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U56 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U57 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U58 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U59 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U60 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U61 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U62 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U63 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U64 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U65 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U66 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U67 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U68 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U69 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U70 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U71 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U72 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U73 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U74 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U75 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U76 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U77 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U78 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U79 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U80 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U81 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U82 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U83 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U84 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U85 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U86 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U87 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U88 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U89 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U90 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U91 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U92 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U93 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U94 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U95 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U96 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U97 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U98 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U99 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U100 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U101 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U102 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U103 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U104 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U105 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U106 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U107 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U108 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U109 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U110 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U111 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U112 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U113 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U114 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U115 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U116 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U117 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U118 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U119 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U120 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U121 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U122 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U123 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U124 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U125 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_15 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n59), .ZN(carry[63]) );
  INV_X1 U3 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U4 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U5 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U6 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U7 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U8 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U9 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U10 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U11 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U12 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U13 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U14 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U15 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U16 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U17 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U18 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U19 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U20 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U21 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U22 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U23 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U24 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U25 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U26 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U27 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U28 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U29 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U30 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U31 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U32 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U33 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U34 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U35 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U36 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U37 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U38 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U39 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U40 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U41 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U42 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U43 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U44 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U45 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U46 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U47 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U48 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U49 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U50 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U51 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U52 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U53 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U54 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U55 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U56 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U57 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U58 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U59 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U60 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U61 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U62 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U63 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U64 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U65 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U66 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U67 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U68 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U69 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U70 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U71 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U72 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U73 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U74 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U75 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U76 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U77 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U78 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U79 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U80 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U81 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U82 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U83 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U84 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U85 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U86 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U87 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U88 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U89 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U90 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U91 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U92 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U93 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U94 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U95 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U96 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  AOI22_X1 U97 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U98 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U99 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U100 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U101 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U102 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U103 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U104 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U105 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U106 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U107 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U108 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U109 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U110 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U111 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U112 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U113 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U114 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U115 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U116 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U117 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U118 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U119 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U120 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U121 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U122 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U123 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U124 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U125 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_16 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  XOR2_X1 U2 ( .A(c[10]), .B(n129), .Z(result[10]) );
  INV_X1 U3 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U4 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U5 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U6 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U7 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U8 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U9 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U10 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U11 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U12 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U13 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U14 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U15 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U16 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U17 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U18 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U19 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U20 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U21 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U22 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U23 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U24 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U25 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U26 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U27 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U28 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U29 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U30 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U31 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U32 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U33 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U34 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U35 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U36 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U37 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U38 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U39 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U40 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U41 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U42 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U43 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U44 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U45 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U46 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U47 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U48 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U49 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U50 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U51 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U52 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U53 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U54 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U55 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U56 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U57 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U58 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U59 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U60 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U61 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U62 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U63 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U64 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U65 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U66 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U67 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U68 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U69 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U70 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U71 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U72 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U73 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U74 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U75 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U76 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U77 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U78 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U79 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U80 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U81 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U82 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U83 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U84 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U85 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U86 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U87 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U88 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U89 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U90 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U91 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U92 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U93 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U94 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U95 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U96 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U97 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U98 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U99 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U100 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U101 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U102 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U103 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U104 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U105 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U106 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U107 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U108 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U109 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U110 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U111 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U112 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U113 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U114 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U115 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U116 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U117 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U118 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U119 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U120 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U121 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U122 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U123 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U124 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U125 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U126 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U127 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U191 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_17 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n207), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n206), .Z(result[8]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n204), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n203), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n203) );
  XOR2_X1 U134 ( .A(c[62]), .B(n202), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n201), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n200), .Z(result[60]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n198), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n197), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n196), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n195), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n194), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n193), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n192), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n191), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n190), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n189), .Z(result[50]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n187), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n186), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n185), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n184), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n183), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n182), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n181), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n180), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n179), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n178), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n177), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n176), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n175), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n174), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n173), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n172), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n171), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n170), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n169), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n168), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n167), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n166), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n165), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n164), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n163), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n162), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n161), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n160), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n159), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n158), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n157), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n156), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n155), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n154), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n153), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n152), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n151), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n150), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n149), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n148), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n147), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n146), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n145), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n144), .Z(result[0]) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n204) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n202) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n201) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n200) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n198) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n197) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n196) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n195) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n194) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n193) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n192) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n191) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n190) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n189) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n187) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n177) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n186) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n185) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n184) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n183) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n182) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n181) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n180) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n179) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n178) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n176) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n166) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n175) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n174) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n173) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n172) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n171) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n170) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n169) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n168) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n167) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n165) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n155) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n164) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n163) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n162) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n161) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n160) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n159) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n158) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n157) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n156) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n154) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n144) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n153) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n152) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n151) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n150) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n149) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n148) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n147) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n146) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n145) );
  INV_X1 U2 ( .A(c[4]), .ZN(n6) );
  INV_X1 U3 ( .A(c[5]), .ZN(n1) );
  INV_X1 U4 ( .A(c[7]), .ZN(n7) );
  INV_X1 U5 ( .A(a[4]), .ZN(n3) );
  INV_X1 U6 ( .A(a[5]), .ZN(n5) );
  INV_X1 U7 ( .A(a[8]), .ZN(n2) );
  INV_X1 U8 ( .A(a[9]), .ZN(n4) );
  XNOR2_X1 U9 ( .A(n199), .B(n1), .ZN(result[5]) );
  XNOR2_X1 U10 ( .A(n2), .B(b[8]), .ZN(n206) );
  XNOR2_X1 U11 ( .A(n3), .B(b[4]), .ZN(n188) );
  XNOR2_X1 U12 ( .A(n4), .B(b[9]), .ZN(n207) );
  XNOR2_X1 U13 ( .A(b[5]), .B(n5), .ZN(n199) );
  XNOR2_X1 U14 ( .A(n6), .B(n188), .ZN(result[4]) );
  XNOR2_X1 U15 ( .A(n205), .B(n7), .ZN(result[7]) );
  INV_X1 U16 ( .A(n58), .ZN(carry[55]) );
  AOI22_X1 U17 ( .A1(b[54]), .A2(a[54]), .B1(n193), .B2(c[54]), .ZN(n58) );
  INV_X1 U18 ( .A(n139), .ZN(carry[63]) );
  AOI22_X1 U19 ( .A1(b[62]), .A2(a[62]), .B1(n202), .B2(c[62]), .ZN(n139) );
  INV_X1 U20 ( .A(n59), .ZN(carry[56]) );
  AOI22_X1 U21 ( .A1(b[55]), .A2(a[55]), .B1(n194), .B2(c[55]), .ZN(n59) );
  INV_X1 U22 ( .A(n60), .ZN(carry[57]) );
  AOI22_X1 U23 ( .A1(b[56]), .A2(a[56]), .B1(n195), .B2(c[56]), .ZN(n60) );
  INV_X1 U24 ( .A(n61), .ZN(carry[58]) );
  AOI22_X1 U25 ( .A1(b[57]), .A2(a[57]), .B1(n196), .B2(c[57]), .ZN(n61) );
  INV_X1 U26 ( .A(n62), .ZN(carry[59]) );
  AOI22_X1 U27 ( .A1(b[58]), .A2(a[58]), .B1(n197), .B2(c[58]), .ZN(n62) );
  INV_X1 U28 ( .A(n136), .ZN(carry[60]) );
  AOI22_X1 U29 ( .A1(b[59]), .A2(a[59]), .B1(n198), .B2(c[59]), .ZN(n136) );
  INV_X1 U30 ( .A(n137), .ZN(carry[61]) );
  AOI22_X1 U31 ( .A1(b[60]), .A2(a[60]), .B1(n200), .B2(c[60]), .ZN(n137) );
  INV_X1 U32 ( .A(n138), .ZN(carry[62]) );
  AOI22_X1 U33 ( .A1(b[61]), .A2(a[61]), .B1(n201), .B2(c[61]), .ZN(n138) );
  INV_X1 U34 ( .A(n21), .ZN(carry[21]) );
  AOI22_X1 U35 ( .A1(b[20]), .A2(a[20]), .B1(n156), .B2(c[20]), .ZN(n21) );
  INV_X1 U36 ( .A(n22), .ZN(carry[22]) );
  AOI22_X1 U37 ( .A1(b[21]), .A2(a[21]), .B1(n157), .B2(c[21]), .ZN(n22) );
  INV_X1 U38 ( .A(n25), .ZN(carry[25]) );
  AOI22_X1 U39 ( .A1(b[24]), .A2(a[24]), .B1(n160), .B2(c[24]), .ZN(n25) );
  INV_X1 U40 ( .A(n26), .ZN(carry[26]) );
  AOI22_X1 U41 ( .A1(b[25]), .A2(a[25]), .B1(n161), .B2(c[25]), .ZN(n26) );
  INV_X1 U42 ( .A(n27), .ZN(carry[27]) );
  AOI22_X1 U43 ( .A1(b[26]), .A2(a[26]), .B1(n162), .B2(c[26]), .ZN(n27) );
  INV_X1 U44 ( .A(n28), .ZN(carry[28]) );
  AOI22_X1 U45 ( .A1(b[27]), .A2(a[27]), .B1(n163), .B2(c[27]), .ZN(n28) );
  INV_X1 U46 ( .A(n29), .ZN(carry[29]) );
  AOI22_X1 U47 ( .A1(b[28]), .A2(a[28]), .B1(n164), .B2(c[28]), .ZN(n29) );
  INV_X1 U48 ( .A(n31), .ZN(carry[30]) );
  AOI22_X1 U49 ( .A1(b[29]), .A2(a[29]), .B1(n165), .B2(c[29]), .ZN(n31) );
  INV_X1 U50 ( .A(a[7]), .ZN(n8) );
  INV_X1 U51 ( .A(n23), .ZN(carry[23]) );
  AOI22_X1 U52 ( .A1(b[22]), .A2(a[22]), .B1(n158), .B2(c[22]), .ZN(n23) );
  INV_X1 U53 ( .A(n24), .ZN(carry[24]) );
  AOI22_X1 U54 ( .A1(b[23]), .A2(a[23]), .B1(n159), .B2(c[23]), .ZN(n24) );
  INV_X1 U55 ( .A(n40), .ZN(carry[39]) );
  AOI22_X1 U56 ( .A1(b[38]), .A2(a[38]), .B1(n175), .B2(c[38]), .ZN(n40) );
  INV_X1 U57 ( .A(n42), .ZN(carry[40]) );
  AOI22_X1 U58 ( .A1(b[39]), .A2(a[39]), .B1(n176), .B2(c[39]), .ZN(n42) );
  INV_X1 U59 ( .A(n43), .ZN(carry[41]) );
  AOI22_X1 U60 ( .A1(b[40]), .A2(a[40]), .B1(n178), .B2(c[40]), .ZN(n43) );
  INV_X1 U61 ( .A(n44), .ZN(carry[42]) );
  AOI22_X1 U62 ( .A1(b[41]), .A2(a[41]), .B1(n179), .B2(c[41]), .ZN(n44) );
  INV_X1 U63 ( .A(n33), .ZN(carry[32]) );
  AOI22_X1 U64 ( .A1(b[31]), .A2(a[31]), .B1(n168), .B2(c[31]), .ZN(n33) );
  INV_X1 U65 ( .A(n34), .ZN(carry[33]) );
  AOI22_X1 U66 ( .A1(b[32]), .A2(a[32]), .B1(n169), .B2(c[32]), .ZN(n34) );
  INV_X1 U67 ( .A(n35), .ZN(carry[34]) );
  AOI22_X1 U68 ( .A1(b[33]), .A2(a[33]), .B1(n170), .B2(c[33]), .ZN(n35) );
  INV_X1 U69 ( .A(n36), .ZN(carry[35]) );
  AOI22_X1 U70 ( .A1(b[34]), .A2(a[34]), .B1(n171), .B2(c[34]), .ZN(n36) );
  INV_X1 U71 ( .A(n37), .ZN(carry[36]) );
  AOI22_X1 U72 ( .A1(b[35]), .A2(a[35]), .B1(n172), .B2(c[35]), .ZN(n37) );
  INV_X1 U73 ( .A(n38), .ZN(carry[37]) );
  AOI22_X1 U74 ( .A1(b[36]), .A2(a[36]), .B1(n173), .B2(c[36]), .ZN(n38) );
  INV_X1 U75 ( .A(n39), .ZN(carry[38]) );
  AOI22_X1 U76 ( .A1(b[37]), .A2(a[37]), .B1(n174), .B2(c[37]), .ZN(n39) );
  INV_X1 U77 ( .A(n32), .ZN(carry[31]) );
  AOI22_X1 U78 ( .A1(b[30]), .A2(a[30]), .B1(n167), .B2(c[30]), .ZN(n32) );
  INV_X1 U79 ( .A(n49), .ZN(carry[47]) );
  AOI22_X1 U80 ( .A1(b[46]), .A2(a[46]), .B1(n184), .B2(c[46]), .ZN(n49) );
  INV_X1 U81 ( .A(n51), .ZN(carry[49]) );
  AOI22_X1 U82 ( .A1(b[48]), .A2(a[48]), .B1(n186), .B2(c[48]), .ZN(n51) );
  INV_X1 U83 ( .A(n54), .ZN(carry[51]) );
  AOI22_X1 U84 ( .A1(b[50]), .A2(a[50]), .B1(n189), .B2(c[50]), .ZN(n54) );
  INV_X1 U85 ( .A(n55), .ZN(carry[52]) );
  AOI22_X1 U86 ( .A1(b[51]), .A2(a[51]), .B1(n190), .B2(c[51]), .ZN(n55) );
  INV_X1 U87 ( .A(n57), .ZN(carry[54]) );
  AOI22_X1 U88 ( .A1(b[53]), .A2(a[53]), .B1(n192), .B2(c[53]), .ZN(n57) );
  INV_X1 U89 ( .A(n45), .ZN(carry[43]) );
  AOI22_X1 U90 ( .A1(b[42]), .A2(a[42]), .B1(n180), .B2(c[42]), .ZN(n45) );
  INV_X1 U91 ( .A(n46), .ZN(carry[44]) );
  AOI22_X1 U92 ( .A1(b[43]), .A2(a[43]), .B1(n181), .B2(c[43]), .ZN(n46) );
  INV_X1 U93 ( .A(n47), .ZN(carry[45]) );
  AOI22_X1 U94 ( .A1(b[44]), .A2(a[44]), .B1(n182), .B2(c[44]), .ZN(n47) );
  INV_X1 U95 ( .A(n48), .ZN(carry[46]) );
  AOI22_X1 U96 ( .A1(b[45]), .A2(a[45]), .B1(n183), .B2(c[45]), .ZN(n48) );
  INV_X1 U97 ( .A(n50), .ZN(carry[48]) );
  AOI22_X1 U98 ( .A1(b[47]), .A2(a[47]), .B1(n185), .B2(c[47]), .ZN(n50) );
  INV_X1 U99 ( .A(n53), .ZN(carry[50]) );
  AOI22_X1 U100 ( .A1(b[49]), .A2(a[49]), .B1(n187), .B2(c[49]), .ZN(n53) );
  INV_X1 U101 ( .A(n56), .ZN(carry[53]) );
  AOI22_X1 U102 ( .A1(b[52]), .A2(a[52]), .B1(n191), .B2(c[52]), .ZN(n56) );
  INV_X1 U103 ( .A(n142), .ZN(carry[8]) );
  INV_X1 U104 ( .A(n143), .ZN(carry[9]) );
  INV_X1 U105 ( .A(n140), .ZN(carry[6]) );
  AOI22_X1 U106 ( .A1(b[5]), .A2(a[5]), .B1(n199), .B2(c[5]), .ZN(n140) );
  INV_X1 U107 ( .A(n141), .ZN(carry[7]) );
  AOI22_X1 U108 ( .A1(b[6]), .A2(a[6]), .B1(n204), .B2(c[6]), .ZN(n141) );
  INV_X1 U109 ( .A(n9), .ZN(carry[10]) );
  AOI22_X1 U110 ( .A1(b[9]), .A2(a[9]), .B1(n207), .B2(c[9]), .ZN(n9) );
  INV_X1 U111 ( .A(n10), .ZN(carry[11]) );
  AOI22_X1 U112 ( .A1(b[10]), .A2(a[10]), .B1(n145), .B2(c[10]), .ZN(n10) );
  INV_X1 U113 ( .A(n11), .ZN(carry[12]) );
  AOI22_X1 U114 ( .A1(b[11]), .A2(a[11]), .B1(n146), .B2(c[11]), .ZN(n11) );
  INV_X1 U115 ( .A(n12), .ZN(carry[13]) );
  AOI22_X1 U116 ( .A1(b[12]), .A2(a[12]), .B1(n147), .B2(c[12]), .ZN(n12) );
  INV_X1 U117 ( .A(n13), .ZN(carry[14]) );
  AOI22_X1 U118 ( .A1(b[13]), .A2(a[13]), .B1(n148), .B2(c[13]), .ZN(n13) );
  INV_X1 U119 ( .A(n14), .ZN(carry[15]) );
  AOI22_X1 U120 ( .A1(b[14]), .A2(a[14]), .B1(n149), .B2(c[14]), .ZN(n14) );
  INV_X1 U121 ( .A(n15), .ZN(carry[16]) );
  AOI22_X1 U122 ( .A1(b[15]), .A2(a[15]), .B1(n150), .B2(c[15]), .ZN(n15) );
  INV_X1 U123 ( .A(n16), .ZN(carry[17]) );
  AOI22_X1 U124 ( .A1(b[16]), .A2(a[16]), .B1(n151), .B2(c[16]), .ZN(n16) );
  INV_X1 U125 ( .A(n17), .ZN(carry[18]) );
  AOI22_X1 U126 ( .A1(b[17]), .A2(a[17]), .B1(n152), .B2(c[17]), .ZN(n17) );
  INV_X1 U127 ( .A(n18), .ZN(carry[19]) );
  AOI22_X1 U130 ( .A1(b[18]), .A2(a[18]), .B1(n153), .B2(c[18]), .ZN(n18) );
  INV_X1 U137 ( .A(n20), .ZN(carry[20]) );
  AOI22_X1 U148 ( .A1(b[19]), .A2(a[19]), .B1(n154), .B2(c[19]), .ZN(n20) );
  INV_X1 U193 ( .A(n30), .ZN(carry[2]) );
  AOI22_X1 U194 ( .A1(b[1]), .A2(a[1]), .B1(n155), .B2(c[1]), .ZN(n30) );
  INV_X1 U196 ( .A(n41), .ZN(carry[3]) );
  AOI22_X1 U201 ( .A1(b[2]), .A2(a[2]), .B1(n166), .B2(c[2]), .ZN(n41) );
  INV_X1 U255 ( .A(n63), .ZN(carry[5]) );
  AOI22_X1 U256 ( .A1(b[4]), .A2(a[4]), .B1(n188), .B2(c[4]), .ZN(n63) );
  INV_X1 U257 ( .A(n52), .ZN(carry[4]) );
  AOI22_X1 U258 ( .A1(b[3]), .A2(a[3]), .B1(n177), .B2(c[3]), .ZN(n52) );
  INV_X1 U259 ( .A(n19), .ZN(carry[1]) );
  AOI22_X1 U260 ( .A1(b[0]), .A2(a[0]), .B1(n144), .B2(c[0]), .ZN(n19) );
  XNOR2_X1 U261 ( .A(b[7]), .B(n8), .ZN(n205) );
  AOI22_X1 U262 ( .A1(b[8]), .A2(a[8]), .B1(n206), .B2(c[8]), .ZN(n143) );
  AOI22_X1 U263 ( .A1(b[7]), .A2(a[7]), .B1(n205), .B2(c[7]), .ZN(n142) );
endmodule


module BWAdder_18 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n235), .Z(result[9]) );
  XOR2_X1 U131 ( .A(n232), .B(c[6]), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n231), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n231) );
  XOR2_X1 U134 ( .A(c[62]), .B(n230), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n229), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n228), .Z(result[60]) );
  XOR2_X1 U137 ( .A(n227), .B(c[5]), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n226), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n225), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n224), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n223), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n222), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n221), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n220), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n219), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n218), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n217), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n216), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n215), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n214), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n213), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n212), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n211), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n210), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n209), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n208), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n207), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n206), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n205), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n204), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n203), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n202), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n201), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n200), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n199), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n198), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n197), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n196), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n195), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n194), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n193), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n192), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n191), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n190), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n189), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n188), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n187), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n186), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n185), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n184), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n183), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n182), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n181), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n180), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n179), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n178), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n177), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n176), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n175), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n174), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n173), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n172), .Z(result[0]) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n230) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n229) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n228) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n226) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n225) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n224) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n223) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n222) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n221) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n220) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n219) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n218) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n217) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n215) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n214) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n213) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n212) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n211) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n210) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n209) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n208) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n207) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n206) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n204) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n194) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n203) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n202) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n201) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n200) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n199) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n198) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n197) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n196) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n195) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n193) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n183) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n192) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n191) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n190) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n189) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n188) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n187) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n186) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n185) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n184) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n182) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n172) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n181) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n180) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n179) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n178) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n177) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n176) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n175) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n174) );
  INV_X1 U2 ( .A(b[10]), .ZN(n3) );
  INV_X1 U3 ( .A(b[3]), .ZN(n13) );
  INV_X1 U4 ( .A(b[4]), .ZN(n7) );
  INV_X1 U5 ( .A(b[5]), .ZN(n19) );
  INV_X1 U6 ( .A(b[6]), .ZN(n18) );
  INV_X1 U7 ( .A(b[9]), .ZN(n12) );
  CLKBUF_X1 U8 ( .A(a[6]), .Z(n1) );
  XOR2_X1 U9 ( .A(a[8]), .B(n21), .Z(n2) );
  INV_X1 U10 ( .A(b[8]), .ZN(n21) );
  XNOR2_X1 U11 ( .A(a[10]), .B(n3), .ZN(n173) );
  NAND2_X1 U12 ( .A1(n234), .A2(n4), .ZN(n5) );
  NAND2_X1 U13 ( .A1(n2), .A2(c[8]), .ZN(n6) );
  NAND2_X1 U14 ( .A1(n6), .A2(n5), .ZN(result[8]) );
  INV_X1 U15 ( .A(c[8]), .ZN(n4) );
  XNOR2_X1 U16 ( .A(a[4]), .B(n7), .ZN(n216) );
  XOR2_X1 U17 ( .A(a[7]), .B(n20), .Z(n8) );
  INV_X1 U18 ( .A(b[7]), .ZN(n20) );
  CLKBUF_X1 U19 ( .A(a[4]), .Z(n9) );
  CLKBUF_X1 U20 ( .A(n234), .Z(n10) );
  CLKBUF_X1 U21 ( .A(a[5]), .Z(n11) );
  XNOR2_X1 U22 ( .A(a[9]), .B(n12), .ZN(n235) );
  XNOR2_X1 U23 ( .A(a[3]), .B(n13), .ZN(n205) );
  CLKBUF_X1 U24 ( .A(n232), .Z(n14) );
  NAND2_X1 U25 ( .A1(n8), .A2(c[7]), .ZN(n16) );
  NAND2_X1 U26 ( .A1(n15), .A2(n233), .ZN(n17) );
  NAND2_X1 U27 ( .A1(n17), .A2(n16), .ZN(result[7]) );
  INV_X1 U28 ( .A(c[7]), .ZN(n15) );
  XNOR2_X1 U29 ( .A(a[6]), .B(n18), .ZN(n232) );
  XNOR2_X1 U30 ( .A(a[5]), .B(n19), .ZN(n227) );
  XNOR2_X1 U31 ( .A(a[7]), .B(n20), .ZN(n233) );
  XNOR2_X1 U32 ( .A(a[8]), .B(n21), .ZN(n234) );
  INV_X1 U33 ( .A(n157), .ZN(carry[54]) );
  AOI22_X1 U34 ( .A1(b[53]), .A2(a[53]), .B1(n220), .B2(c[53]), .ZN(n157) );
  INV_X1 U35 ( .A(n158), .ZN(carry[55]) );
  AOI22_X1 U36 ( .A1(b[54]), .A2(a[54]), .B1(n221), .B2(c[54]), .ZN(n158) );
  INV_X1 U37 ( .A(n159), .ZN(carry[56]) );
  AOI22_X1 U38 ( .A1(b[55]), .A2(a[55]), .B1(n222), .B2(c[55]), .ZN(n159) );
  INV_X1 U39 ( .A(n160), .ZN(carry[57]) );
  AOI22_X1 U40 ( .A1(b[56]), .A2(a[56]), .B1(n223), .B2(c[56]), .ZN(n160) );
  INV_X1 U41 ( .A(n161), .ZN(carry[58]) );
  AOI22_X1 U42 ( .A1(b[57]), .A2(a[57]), .B1(n224), .B2(c[57]), .ZN(n161) );
  INV_X1 U43 ( .A(n162), .ZN(carry[59]) );
  AOI22_X1 U44 ( .A1(b[58]), .A2(a[58]), .B1(n225), .B2(c[58]), .ZN(n162) );
  INV_X1 U45 ( .A(n164), .ZN(carry[60]) );
  AOI22_X1 U46 ( .A1(b[59]), .A2(a[59]), .B1(n226), .B2(c[59]), .ZN(n164) );
  INV_X1 U47 ( .A(n165), .ZN(carry[61]) );
  AOI22_X1 U48 ( .A1(b[60]), .A2(a[60]), .B1(n228), .B2(c[60]), .ZN(n165) );
  INV_X1 U49 ( .A(n166), .ZN(carry[62]) );
  AOI22_X1 U50 ( .A1(b[61]), .A2(a[61]), .B1(n229), .B2(c[61]), .ZN(n166) );
  INV_X1 U51 ( .A(n167), .ZN(carry[63]) );
  AOI22_X1 U52 ( .A1(b[62]), .A2(a[62]), .B1(n230), .B2(c[62]), .ZN(n167) );
  INV_X1 U53 ( .A(n163), .ZN(carry[5]) );
  INV_X1 U54 ( .A(n152), .ZN(carry[4]) );
  INV_X1 U55 ( .A(n168), .ZN(carry[6]) );
  INV_X1 U56 ( .A(n170), .ZN(carry[8]) );
  INV_X1 U57 ( .A(n171), .ZN(carry[9]) );
  INV_X1 U58 ( .A(n169), .ZN(carry[7]) );
  INV_X1 U59 ( .A(n24), .ZN(carry[11]) );
  INV_X1 U60 ( .A(n23), .ZN(carry[10]) );
  INV_X1 U61 ( .A(n42), .ZN(carry[28]) );
  AOI22_X1 U62 ( .A1(b[27]), .A2(a[27]), .B1(n191), .B2(c[27]), .ZN(n42) );
  INV_X1 U63 ( .A(n43), .ZN(carry[29]) );
  AOI22_X1 U64 ( .A1(b[28]), .A2(a[28]), .B1(n192), .B2(c[28]), .ZN(n43) );
  INV_X1 U65 ( .A(n45), .ZN(carry[30]) );
  AOI22_X1 U66 ( .A1(b[29]), .A2(a[29]), .B1(n193), .B2(c[29]), .ZN(n45) );
  INV_X1 U67 ( .A(n32), .ZN(carry[19]) );
  AOI22_X1 U68 ( .A1(b[18]), .A2(a[18]), .B1(n181), .B2(c[18]), .ZN(n32) );
  INV_X1 U69 ( .A(n35), .ZN(carry[21]) );
  AOI22_X1 U70 ( .A1(b[20]), .A2(a[20]), .B1(n184), .B2(c[20]), .ZN(n35) );
  INV_X1 U71 ( .A(n30), .ZN(carry[17]) );
  AOI22_X1 U72 ( .A1(b[16]), .A2(a[16]), .B1(n179), .B2(c[16]), .ZN(n30) );
  INV_X1 U73 ( .A(n34), .ZN(carry[20]) );
  AOI22_X1 U74 ( .A1(b[19]), .A2(a[19]), .B1(n182), .B2(c[19]), .ZN(n34) );
  INV_X1 U75 ( .A(n25), .ZN(carry[12]) );
  AOI22_X1 U76 ( .A1(b[11]), .A2(a[11]), .B1(n174), .B2(c[11]), .ZN(n25) );
  INV_X1 U77 ( .A(n55), .ZN(carry[3]) );
  AOI22_X1 U78 ( .A1(b[2]), .A2(a[2]), .B1(n194), .B2(c[2]), .ZN(n55) );
  INV_X1 U79 ( .A(n26), .ZN(carry[13]) );
  AOI22_X1 U80 ( .A1(b[12]), .A2(a[12]), .B1(n175), .B2(c[12]), .ZN(n26) );
  INV_X1 U81 ( .A(n27), .ZN(carry[14]) );
  AOI22_X1 U82 ( .A1(b[13]), .A2(a[13]), .B1(n176), .B2(c[13]), .ZN(n27) );
  INV_X1 U83 ( .A(n28), .ZN(carry[15]) );
  AOI22_X1 U84 ( .A1(b[14]), .A2(a[14]), .B1(n177), .B2(c[14]), .ZN(n28) );
  INV_X1 U85 ( .A(n31), .ZN(carry[18]) );
  AOI22_X1 U86 ( .A1(b[17]), .A2(a[17]), .B1(n180), .B2(c[17]), .ZN(n31) );
  INV_X1 U87 ( .A(n29), .ZN(carry[16]) );
  AOI22_X1 U88 ( .A1(b[15]), .A2(a[15]), .B1(n178), .B2(c[15]), .ZN(n29) );
  INV_X1 U89 ( .A(n36), .ZN(carry[22]) );
  AOI22_X1 U90 ( .A1(b[21]), .A2(a[21]), .B1(n185), .B2(c[21]), .ZN(n36) );
  INV_X1 U91 ( .A(n37), .ZN(carry[23]) );
  AOI22_X1 U92 ( .A1(b[22]), .A2(a[22]), .B1(n186), .B2(c[22]), .ZN(n37) );
  INV_X1 U93 ( .A(n38), .ZN(carry[24]) );
  AOI22_X1 U94 ( .A1(b[23]), .A2(a[23]), .B1(n187), .B2(c[23]), .ZN(n38) );
  INV_X1 U95 ( .A(n39), .ZN(carry[25]) );
  AOI22_X1 U96 ( .A1(b[24]), .A2(a[24]), .B1(n188), .B2(c[24]), .ZN(n39) );
  INV_X1 U97 ( .A(n40), .ZN(carry[26]) );
  AOI22_X1 U98 ( .A1(b[25]), .A2(a[25]), .B1(n189), .B2(c[25]), .ZN(n40) );
  INV_X1 U99 ( .A(n41), .ZN(carry[27]) );
  AOI22_X1 U100 ( .A1(b[26]), .A2(a[26]), .B1(n190), .B2(c[26]), .ZN(n41) );
  INV_X1 U101 ( .A(n46), .ZN(carry[31]) );
  AOI22_X1 U102 ( .A1(b[30]), .A2(a[30]), .B1(n195), .B2(c[30]), .ZN(n46) );
  INV_X1 U103 ( .A(n47), .ZN(carry[32]) );
  AOI22_X1 U104 ( .A1(b[31]), .A2(a[31]), .B1(n196), .B2(c[31]), .ZN(n47) );
  INV_X1 U105 ( .A(n48), .ZN(carry[33]) );
  AOI22_X1 U106 ( .A1(b[32]), .A2(a[32]), .B1(n197), .B2(c[32]), .ZN(n48) );
  INV_X1 U107 ( .A(n49), .ZN(carry[34]) );
  AOI22_X1 U108 ( .A1(b[33]), .A2(a[33]), .B1(n198), .B2(c[33]), .ZN(n49) );
  INV_X1 U109 ( .A(n50), .ZN(carry[35]) );
  AOI22_X1 U110 ( .A1(b[34]), .A2(a[34]), .B1(n199), .B2(c[34]), .ZN(n50) );
  INV_X1 U111 ( .A(n51), .ZN(carry[36]) );
  AOI22_X1 U112 ( .A1(b[35]), .A2(a[35]), .B1(n200), .B2(c[35]), .ZN(n51) );
  INV_X1 U113 ( .A(n52), .ZN(carry[37]) );
  AOI22_X1 U114 ( .A1(b[36]), .A2(a[36]), .B1(n201), .B2(c[36]), .ZN(n52) );
  INV_X1 U115 ( .A(n53), .ZN(carry[38]) );
  AOI22_X1 U116 ( .A1(b[37]), .A2(a[37]), .B1(n202), .B2(c[37]), .ZN(n53) );
  INV_X1 U117 ( .A(n54), .ZN(carry[39]) );
  AOI22_X1 U118 ( .A1(b[38]), .A2(a[38]), .B1(n203), .B2(c[38]), .ZN(n54) );
  INV_X1 U119 ( .A(n56), .ZN(carry[40]) );
  AOI22_X1 U120 ( .A1(b[39]), .A2(a[39]), .B1(n204), .B2(c[39]), .ZN(n56) );
  INV_X1 U121 ( .A(n57), .ZN(carry[41]) );
  AOI22_X1 U122 ( .A1(b[40]), .A2(a[40]), .B1(n206), .B2(c[40]), .ZN(n57) );
  INV_X1 U123 ( .A(n58), .ZN(carry[42]) );
  AOI22_X1 U124 ( .A1(b[41]), .A2(a[41]), .B1(n207), .B2(c[41]), .ZN(n58) );
  INV_X1 U125 ( .A(n59), .ZN(carry[43]) );
  AOI22_X1 U126 ( .A1(b[42]), .A2(a[42]), .B1(n208), .B2(c[42]), .ZN(n59) );
  INV_X1 U127 ( .A(n61), .ZN(carry[45]) );
  AOI22_X1 U129 ( .A1(b[44]), .A2(a[44]), .B1(n210), .B2(c[44]), .ZN(n61) );
  INV_X1 U130 ( .A(n62), .ZN(carry[46]) );
  AOI22_X1 U193 ( .A1(b[45]), .A2(a[45]), .B1(n211), .B2(c[45]), .ZN(n62) );
  INV_X1 U194 ( .A(n151), .ZN(carry[49]) );
  AOI22_X1 U195 ( .A1(b[48]), .A2(a[48]), .B1(n214), .B2(c[48]), .ZN(n151) );
  INV_X1 U196 ( .A(n60), .ZN(carry[44]) );
  AOI22_X1 U201 ( .A1(b[43]), .A2(a[43]), .B1(n209), .B2(c[43]), .ZN(n60) );
  INV_X1 U212 ( .A(n63), .ZN(carry[47]) );
  AOI22_X1 U254 ( .A1(b[46]), .A2(a[46]), .B1(n212), .B2(c[46]), .ZN(n63) );
  INV_X1 U255 ( .A(n150), .ZN(carry[48]) );
  AOI22_X1 U256 ( .A1(b[47]), .A2(a[47]), .B1(n213), .B2(c[47]), .ZN(n150) );
  INV_X1 U257 ( .A(n153), .ZN(carry[50]) );
  AOI22_X1 U258 ( .A1(b[49]), .A2(a[49]), .B1(n215), .B2(c[49]), .ZN(n153) );
  INV_X1 U259 ( .A(n154), .ZN(carry[51]) );
  AOI22_X1 U260 ( .A1(b[50]), .A2(a[50]), .B1(n217), .B2(c[50]), .ZN(n154) );
  INV_X1 U261 ( .A(n155), .ZN(carry[52]) );
  AOI22_X1 U262 ( .A1(b[51]), .A2(a[51]), .B1(n218), .B2(c[51]), .ZN(n155) );
  INV_X1 U263 ( .A(n156), .ZN(carry[53]) );
  AOI22_X1 U264 ( .A1(b[52]), .A2(a[52]), .B1(n219), .B2(c[52]), .ZN(n156) );
  INV_X1 U265 ( .A(n44), .ZN(carry[2]) );
  AOI22_X1 U266 ( .A1(b[1]), .A2(a[1]), .B1(n183), .B2(c[1]), .ZN(n44) );
  INV_X1 U267 ( .A(n33), .ZN(carry[1]) );
  AOI22_X1 U268 ( .A1(b[0]), .A2(a[0]), .B1(n172), .B2(c[0]), .ZN(n33) );
  AOI22_X1 U269 ( .A1(b[3]), .A2(a[3]), .B1(n205), .B2(c[3]), .ZN(n152) );
  CLKBUF_X1 U270 ( .A(a[8]), .Z(n22) );
  AOI22_X1 U271 ( .A1(b[9]), .A2(a[9]), .B1(n235), .B2(c[9]), .ZN(n23) );
  AOI22_X1 U272 ( .A1(b[4]), .A2(n9), .B1(n216), .B2(c[4]), .ZN(n163) );
  AOI22_X1 U273 ( .A1(b[10]), .A2(a[10]), .B1(n173), .B2(c[10]), .ZN(n24) );
  AOI22_X1 U274 ( .A1(b[8]), .A2(n22), .B1(n10), .B2(c[8]), .ZN(n171) );
  AOI22_X1 U275 ( .A1(b[5]), .A2(n11), .B1(n227), .B2(c[5]), .ZN(n168) );
  AOI22_X1 U276 ( .A1(b[7]), .A2(a[7]), .B1(n233), .B2(c[7]), .ZN(n170) );
  AOI22_X1 U277 ( .A1(b[6]), .A2(n1), .B1(n14), .B2(c[6]), .ZN(n169) );
endmodule


module BWAdder_19 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n59), .ZN(carry[63]) );
  INV_X1 U3 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U4 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U5 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U6 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U7 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U8 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U9 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U10 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  AOI22_X1 U11 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U12 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U13 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U14 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U15 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U16 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U17 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U18 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U19 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U20 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U21 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U22 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U23 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U24 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U25 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U26 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U27 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U28 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U29 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U30 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U31 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U32 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U33 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U34 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U35 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U36 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U37 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U38 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U39 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U40 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U41 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U42 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U43 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U44 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U45 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U46 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U47 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U48 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U49 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U50 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U51 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U52 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U53 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U54 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U55 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U56 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U57 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U58 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U59 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U60 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U61 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U62 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U63 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U64 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U65 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U66 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U67 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U68 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U69 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U70 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U71 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U72 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U73 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U74 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U75 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U76 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U77 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U78 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U79 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U80 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U81 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U82 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U83 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U84 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U85 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U86 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U87 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U88 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U89 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U90 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U91 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U92 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U93 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U94 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U95 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U96 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U97 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U98 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U99 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U100 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U101 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U102 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U103 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U104 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U105 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U106 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U107 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U108 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U109 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U110 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U111 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U112 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U113 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U114 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U115 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U116 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U117 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U118 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U119 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U120 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U121 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U122 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U123 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U124 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U125 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_20 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U3 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U4 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U5 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U6 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U7 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U8 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U9 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U10 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U11 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U12 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U13 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U14 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U15 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U16 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U17 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U18 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U19 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U20 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U21 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U22 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U23 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U24 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U25 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U26 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U27 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U28 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U29 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U30 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U31 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U32 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U33 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U34 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U35 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U36 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U37 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U38 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U39 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U40 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U41 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U42 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U43 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U44 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U45 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U46 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U47 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U48 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U49 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U50 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U51 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U52 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U53 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U54 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U55 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U56 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U57 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U58 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U59 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U60 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U61 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U62 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U63 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U64 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U65 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U66 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U67 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U68 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U69 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U70 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U71 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U72 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U73 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U74 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U75 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U76 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U77 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U78 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U79 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U80 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U81 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U82 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U83 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U84 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U85 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U86 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U87 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U88 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U89 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U90 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U91 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U92 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U93 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U94 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U95 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U96 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U97 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U98 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U99 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U100 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U101 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U102 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U103 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U104 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U105 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U106 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U107 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U108 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U109 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U110 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U111 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U112 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U113 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U114 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U115 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U116 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U117 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U118 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U119 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U120 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U121 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U122 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U123 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U124 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U125 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_21 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U3 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U4 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U5 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U6 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U7 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U8 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U9 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U10 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U11 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U12 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U13 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U14 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U15 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U16 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U17 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U18 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U19 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U20 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U21 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U22 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U23 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U24 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U25 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U26 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U27 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U28 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U29 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U30 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U31 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U32 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U33 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U34 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U35 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U36 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U37 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U38 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U39 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U40 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U41 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U42 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U43 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U44 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U45 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U46 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U47 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U48 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U49 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U50 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U51 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U52 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U53 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U54 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U55 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U56 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U57 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U58 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U59 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U60 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U61 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U62 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U63 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U64 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U65 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U66 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U67 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U68 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U69 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U70 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U71 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U72 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U73 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U74 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U75 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U76 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U77 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U78 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U79 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U80 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U81 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U82 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U83 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U84 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U85 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U86 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U87 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U88 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U89 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U90 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U91 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U92 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U93 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U94 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U95 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U96 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U97 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U98 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U99 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U100 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U101 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U102 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U103 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U104 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U105 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U106 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U107 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U108 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U109 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U110 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U111 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U112 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U113 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U114 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U115 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U116 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U117 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U118 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U119 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U120 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U121 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U122 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U123 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U124 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U125 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_22 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U3 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U4 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U5 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U6 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U7 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U8 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U9 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U10 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U11 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U12 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U13 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U14 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U15 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U16 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U17 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U18 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U19 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U20 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U21 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U22 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U23 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U24 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U25 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U26 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U27 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U28 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U29 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U30 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U31 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U32 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U33 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U34 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U35 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U36 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U37 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U38 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U39 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U40 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U41 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U42 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U43 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U44 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U45 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U46 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U47 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U48 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U49 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U50 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U51 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U52 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U53 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U55 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U57 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U59 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U61 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U62 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U63 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U64 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U65 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U66 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U67 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U68 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U69 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U70 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U71 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U72 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U73 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U74 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U75 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U76 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U77 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U78 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U79 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U80 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U81 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U82 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U83 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U84 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U85 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U86 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U87 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U88 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U89 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U90 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U91 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U92 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U93 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U94 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U95 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U96 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U97 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U98 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U99 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U100 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U101 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U102 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U103 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U104 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U105 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U106 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U107 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U108 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U109 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U110 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U111 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U112 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U113 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U114 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U115 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U116 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U117 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U118 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U119 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U120 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U121 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U122 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U123 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U124 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U125 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_23 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n215), .Z(result[9]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n212), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n211), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n211) );
  XOR2_X1 U134 ( .A(c[62]), .B(n210), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n209), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n208), .Z(result[60]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n206), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n205), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n204), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n203), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n202), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n201), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n200), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n199), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n198), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n197), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n196), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n195), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n194), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n193), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n192), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n191), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n190), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n189), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n188), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n187), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n186), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n185), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n184), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n183), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n182), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n181), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n180), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n179), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n178), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n177), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n176), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n175), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n174), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n173), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n172), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n171), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n170), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n169), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n168), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n167), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n166), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n165), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n164), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n163), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n162), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n161), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n160), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n159), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n158), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n157), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n156), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n155), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n154), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n153), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n152), .Z(result[0]) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n212) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n210) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n209) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n208) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n206) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n205) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n204) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n203) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n202) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n201) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n200) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n199) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n198) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n197) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n195) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n185) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n194) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n193) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n192) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n191) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n190) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n189) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n188) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n187) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n186) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n184) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n174) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n183) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n182) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n181) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n180) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n179) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n178) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n177) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n176) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n175) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n173) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n163) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n172) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n171) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n170) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n169) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n168) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n167) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n166) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n165) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n164) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n162) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n152) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n161) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n160) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n159) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n158) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n157) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n156) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n155) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n154) );
  INV_X1 U2 ( .A(b[8]), .ZN(n9) );
  INV_X1 U3 ( .A(b[7]), .ZN(n11) );
  INV_X1 U4 ( .A(b[5]), .ZN(n8) );
  INV_X1 U5 ( .A(b[9]), .ZN(n7) );
  INV_X1 U6 ( .A(b[4]), .ZN(n10) );
  INV_X1 U7 ( .A(c[8]), .ZN(n5) );
  INV_X1 U8 ( .A(c[7]), .ZN(n12) );
  INV_X1 U9 ( .A(c[5]), .ZN(n6) );
  NAND2_X1 U10 ( .A1(a[10]), .A2(n2), .ZN(n3) );
  NAND2_X1 U11 ( .A1(n1), .A2(b[10]), .ZN(n4) );
  NAND2_X1 U12 ( .A1(n3), .A2(n4), .ZN(n153) );
  INV_X1 U13 ( .A(a[10]), .ZN(n1) );
  INV_X1 U14 ( .A(b[10]), .ZN(n2) );
  XNOR2_X1 U15 ( .A(n5), .B(n214), .ZN(result[8]) );
  XNOR2_X1 U16 ( .A(n207), .B(n6), .ZN(result[5]) );
  XNOR2_X1 U17 ( .A(a[9]), .B(n7), .ZN(n215) );
  XNOR2_X1 U18 ( .A(a[5]), .B(n8), .ZN(n207) );
  XNOR2_X1 U19 ( .A(a[8]), .B(n9), .ZN(n214) );
  XNOR2_X1 U20 ( .A(a[4]), .B(n10), .ZN(n196) );
  XNOR2_X1 U21 ( .A(a[7]), .B(n11), .ZN(n213) );
  XNOR2_X1 U22 ( .A(n213), .B(n12), .ZN(result[7]) );
  INV_X1 U23 ( .A(n32), .ZN(carry[28]) );
  AOI22_X1 U24 ( .A1(b[27]), .A2(a[27]), .B1(n171), .B2(c[27]), .ZN(n32) );
  INV_X1 U25 ( .A(n33), .ZN(carry[29]) );
  AOI22_X1 U26 ( .A1(b[28]), .A2(a[28]), .B1(n172), .B2(c[28]), .ZN(n33) );
  INV_X1 U27 ( .A(n35), .ZN(carry[30]) );
  AOI22_X1 U28 ( .A1(b[29]), .A2(a[29]), .B1(n173), .B2(c[29]), .ZN(n35) );
  INV_X1 U29 ( .A(n36), .ZN(carry[31]) );
  AOI22_X1 U30 ( .A1(b[30]), .A2(a[30]), .B1(n175), .B2(c[30]), .ZN(n36) );
  INV_X1 U31 ( .A(n37), .ZN(carry[32]) );
  AOI22_X1 U32 ( .A1(b[31]), .A2(a[31]), .B1(n176), .B2(c[31]), .ZN(n37) );
  INV_X1 U33 ( .A(n39), .ZN(carry[34]) );
  AOI22_X1 U34 ( .A1(b[33]), .A2(a[33]), .B1(n178), .B2(c[33]), .ZN(n39) );
  INV_X1 U35 ( .A(n38), .ZN(carry[33]) );
  AOI22_X1 U36 ( .A1(b[32]), .A2(a[32]), .B1(n177), .B2(c[32]), .ZN(n38) );
  INV_X1 U37 ( .A(n40), .ZN(carry[35]) );
  AOI22_X1 U38 ( .A1(b[34]), .A2(a[34]), .B1(n179), .B2(c[34]), .ZN(n40) );
  INV_X1 U39 ( .A(n41), .ZN(carry[36]) );
  AOI22_X1 U40 ( .A1(b[35]), .A2(a[35]), .B1(n180), .B2(c[35]), .ZN(n41) );
  INV_X1 U41 ( .A(n42), .ZN(carry[37]) );
  AOI22_X1 U42 ( .A1(b[36]), .A2(a[36]), .B1(n181), .B2(c[36]), .ZN(n42) );
  INV_X1 U43 ( .A(n43), .ZN(carry[38]) );
  AOI22_X1 U44 ( .A1(b[37]), .A2(a[37]), .B1(n182), .B2(c[37]), .ZN(n43) );
  INV_X1 U45 ( .A(n44), .ZN(carry[39]) );
  AOI22_X1 U46 ( .A1(b[38]), .A2(a[38]), .B1(n183), .B2(c[38]), .ZN(n44) );
  INV_X1 U47 ( .A(n46), .ZN(carry[40]) );
  AOI22_X1 U48 ( .A1(b[39]), .A2(a[39]), .B1(n184), .B2(c[39]), .ZN(n46) );
  INV_X1 U49 ( .A(n47), .ZN(carry[41]) );
  AOI22_X1 U50 ( .A1(b[40]), .A2(a[40]), .B1(n186), .B2(c[40]), .ZN(n47) );
  INV_X1 U51 ( .A(n48), .ZN(carry[42]) );
  AOI22_X1 U52 ( .A1(b[41]), .A2(a[41]), .B1(n187), .B2(c[41]), .ZN(n48) );
  INV_X1 U53 ( .A(n49), .ZN(carry[43]) );
  AOI22_X1 U54 ( .A1(b[42]), .A2(a[42]), .B1(n188), .B2(c[42]), .ZN(n49) );
  INV_X1 U55 ( .A(n50), .ZN(carry[44]) );
  AOI22_X1 U56 ( .A1(b[43]), .A2(a[43]), .B1(n189), .B2(c[43]), .ZN(n50) );
  INV_X1 U57 ( .A(n51), .ZN(carry[45]) );
  AOI22_X1 U58 ( .A1(b[44]), .A2(a[44]), .B1(n190), .B2(c[44]), .ZN(n51) );
  INV_X1 U59 ( .A(n52), .ZN(carry[46]) );
  AOI22_X1 U60 ( .A1(b[45]), .A2(a[45]), .B1(n191), .B2(c[45]), .ZN(n52) );
  INV_X1 U61 ( .A(n53), .ZN(carry[47]) );
  AOI22_X1 U62 ( .A1(b[46]), .A2(a[46]), .B1(n192), .B2(c[46]), .ZN(n53) );
  INV_X1 U63 ( .A(n54), .ZN(carry[48]) );
  AOI22_X1 U64 ( .A1(b[47]), .A2(a[47]), .B1(n193), .B2(c[47]), .ZN(n54) );
  INV_X1 U65 ( .A(n55), .ZN(carry[49]) );
  AOI22_X1 U66 ( .A1(b[48]), .A2(a[48]), .B1(n194), .B2(c[48]), .ZN(n55) );
  INV_X1 U67 ( .A(n57), .ZN(carry[50]) );
  AOI22_X1 U68 ( .A1(b[49]), .A2(a[49]), .B1(n195), .B2(c[49]), .ZN(n57) );
  INV_X1 U69 ( .A(n58), .ZN(carry[51]) );
  AOI22_X1 U70 ( .A1(b[50]), .A2(a[50]), .B1(n197), .B2(c[50]), .ZN(n58) );
  INV_X1 U71 ( .A(n59), .ZN(carry[52]) );
  AOI22_X1 U72 ( .A1(b[51]), .A2(a[51]), .B1(n198), .B2(c[51]), .ZN(n59) );
  INV_X1 U73 ( .A(n60), .ZN(carry[53]) );
  AOI22_X1 U74 ( .A1(b[52]), .A2(a[52]), .B1(n199), .B2(c[52]), .ZN(n60) );
  INV_X1 U75 ( .A(n61), .ZN(carry[54]) );
  AOI22_X1 U76 ( .A1(b[53]), .A2(a[53]), .B1(n200), .B2(c[53]), .ZN(n61) );
  INV_X1 U77 ( .A(n62), .ZN(carry[55]) );
  AOI22_X1 U78 ( .A1(b[54]), .A2(a[54]), .B1(n201), .B2(c[54]), .ZN(n62) );
  INV_X1 U79 ( .A(n63), .ZN(carry[56]) );
  AOI22_X1 U80 ( .A1(b[55]), .A2(a[55]), .B1(n202), .B2(c[55]), .ZN(n63) );
  INV_X1 U81 ( .A(n147), .ZN(carry[63]) );
  INV_X1 U82 ( .A(n140), .ZN(carry[57]) );
  AOI22_X1 U83 ( .A1(b[56]), .A2(a[56]), .B1(n203), .B2(c[56]), .ZN(n140) );
  INV_X1 U84 ( .A(n141), .ZN(carry[58]) );
  AOI22_X1 U85 ( .A1(b[57]), .A2(a[57]), .B1(n204), .B2(c[57]), .ZN(n141) );
  INV_X1 U86 ( .A(n142), .ZN(carry[59]) );
  AOI22_X1 U87 ( .A1(b[58]), .A2(a[58]), .B1(n205), .B2(c[58]), .ZN(n142) );
  AOI22_X1 U88 ( .A1(b[62]), .A2(a[62]), .B1(n210), .B2(c[62]), .ZN(n147) );
  INV_X1 U89 ( .A(n144), .ZN(carry[60]) );
  AOI22_X1 U90 ( .A1(b[59]), .A2(a[59]), .B1(n206), .B2(c[59]), .ZN(n144) );
  INV_X1 U91 ( .A(n145), .ZN(carry[61]) );
  AOI22_X1 U92 ( .A1(b[60]), .A2(a[60]), .B1(n208), .B2(c[60]), .ZN(n145) );
  INV_X1 U93 ( .A(n146), .ZN(carry[62]) );
  AOI22_X1 U94 ( .A1(b[61]), .A2(a[61]), .B1(n209), .B2(c[61]), .ZN(n146) );
  INV_X1 U95 ( .A(n27), .ZN(carry[23]) );
  AOI22_X1 U96 ( .A1(b[22]), .A2(a[22]), .B1(n166), .B2(c[22]), .ZN(n27) );
  INV_X1 U97 ( .A(n28), .ZN(carry[24]) );
  AOI22_X1 U98 ( .A1(b[23]), .A2(a[23]), .B1(n167), .B2(c[23]), .ZN(n28) );
  INV_X1 U99 ( .A(n29), .ZN(carry[25]) );
  AOI22_X1 U100 ( .A1(b[24]), .A2(a[24]), .B1(n168), .B2(c[24]), .ZN(n29) );
  INV_X1 U101 ( .A(n30), .ZN(carry[26]) );
  AOI22_X1 U102 ( .A1(b[25]), .A2(a[25]), .B1(n169), .B2(c[25]), .ZN(n30) );
  INV_X1 U103 ( .A(n31), .ZN(carry[27]) );
  AOI22_X1 U104 ( .A1(b[26]), .A2(a[26]), .B1(n170), .B2(c[26]), .ZN(n31) );
  INV_X1 U105 ( .A(n25), .ZN(carry[21]) );
  AOI22_X1 U106 ( .A1(b[20]), .A2(a[20]), .B1(n164), .B2(c[20]), .ZN(n25) );
  INV_X1 U107 ( .A(n26), .ZN(carry[22]) );
  AOI22_X1 U108 ( .A1(b[21]), .A2(a[21]), .B1(n165), .B2(c[21]), .ZN(n26) );
  INV_X1 U109 ( .A(n21), .ZN(carry[18]) );
  AOI22_X1 U110 ( .A1(b[17]), .A2(a[17]), .B1(n160), .B2(c[17]), .ZN(n21) );
  INV_X1 U111 ( .A(n24), .ZN(carry[20]) );
  AOI22_X1 U112 ( .A1(b[19]), .A2(a[19]), .B1(n162), .B2(c[19]), .ZN(n24) );
  INV_X1 U113 ( .A(n22), .ZN(carry[19]) );
  AOI22_X1 U114 ( .A1(b[18]), .A2(a[18]), .B1(n161), .B2(c[18]), .ZN(n22) );
  INV_X1 U115 ( .A(n20), .ZN(carry[17]) );
  AOI22_X1 U116 ( .A1(b[16]), .A2(a[16]), .B1(n159), .B2(c[16]), .ZN(n20) );
  INV_X1 U117 ( .A(n19), .ZN(carry[16]) );
  AOI22_X1 U118 ( .A1(b[15]), .A2(a[15]), .B1(n158), .B2(c[15]), .ZN(n19) );
  INV_X1 U119 ( .A(n17), .ZN(carry[14]) );
  AOI22_X1 U120 ( .A1(b[13]), .A2(a[13]), .B1(n156), .B2(c[13]), .ZN(n17) );
  INV_X1 U121 ( .A(n18), .ZN(carry[15]) );
  AOI22_X1 U122 ( .A1(b[14]), .A2(a[14]), .B1(n157), .B2(c[14]), .ZN(n18) );
  INV_X1 U123 ( .A(n150), .ZN(carry[8]) );
  INV_X1 U124 ( .A(n151), .ZN(carry[9]) );
  INV_X1 U125 ( .A(n143), .ZN(carry[5]) );
  AOI22_X1 U126 ( .A1(b[4]), .A2(a[4]), .B1(n196), .B2(c[4]), .ZN(n143) );
  INV_X1 U127 ( .A(n148), .ZN(carry[6]) );
  AOI22_X1 U129 ( .A1(b[5]), .A2(a[5]), .B1(n207), .B2(c[5]), .ZN(n148) );
  INV_X1 U130 ( .A(n149), .ZN(carry[7]) );
  AOI22_X1 U137 ( .A1(b[6]), .A2(a[6]), .B1(n212), .B2(c[6]), .ZN(n149) );
  INV_X1 U193 ( .A(n13), .ZN(carry[10]) );
  AOI22_X1 U194 ( .A1(b[9]), .A2(a[9]), .B1(n215), .B2(c[9]), .ZN(n13) );
  INV_X1 U196 ( .A(n14), .ZN(carry[11]) );
  AOI22_X1 U201 ( .A1(b[10]), .A2(a[10]), .B1(n153), .B2(c[10]), .ZN(n14) );
  INV_X1 U254 ( .A(n15), .ZN(carry[12]) );
  AOI22_X1 U255 ( .A1(b[11]), .A2(a[11]), .B1(n154), .B2(c[11]), .ZN(n15) );
  INV_X1 U256 ( .A(n16), .ZN(carry[13]) );
  AOI22_X1 U257 ( .A1(b[12]), .A2(a[12]), .B1(n155), .B2(c[12]), .ZN(n16) );
  INV_X1 U258 ( .A(n34), .ZN(carry[2]) );
  AOI22_X1 U259 ( .A1(b[1]), .A2(a[1]), .B1(n163), .B2(c[1]), .ZN(n34) );
  INV_X1 U260 ( .A(n45), .ZN(carry[3]) );
  AOI22_X1 U261 ( .A1(b[2]), .A2(a[2]), .B1(n174), .B2(c[2]), .ZN(n45) );
  INV_X1 U262 ( .A(n56), .ZN(carry[4]) );
  AOI22_X1 U263 ( .A1(b[3]), .A2(a[3]), .B1(n185), .B2(c[3]), .ZN(n56) );
  INV_X1 U264 ( .A(n23), .ZN(carry[1]) );
  AOI22_X1 U265 ( .A1(b[0]), .A2(a[0]), .B1(n152), .B2(c[0]), .ZN(n23) );
  AOI22_X1 U266 ( .A1(b[8]), .A2(a[8]), .B1(n214), .B2(c[8]), .ZN(n151) );
  AOI22_X1 U267 ( .A1(b[7]), .A2(a[7]), .B1(n213), .B2(c[7]), .ZN(n150) );
endmodule


module BWAdder_24 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U3 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U4 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U5 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U6 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U7 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U8 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U9 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U10 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U11 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U12 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U13 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U14 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U15 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U16 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U17 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U18 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U19 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U20 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U21 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U22 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U23 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U24 ( .A(n59), .ZN(carry[63]) );
  INV_X1 U25 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U26 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U27 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U28 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U29 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U30 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U31 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U32 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U33 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U34 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U35 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U36 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  AOI22_X1 U37 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U38 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U39 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U40 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U41 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U42 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U43 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U44 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U45 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U46 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U47 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U48 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U49 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U50 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U51 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U52 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U53 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U54 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U55 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U56 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U57 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U58 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U59 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U60 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U61 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U62 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U63 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U64 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U65 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U66 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U67 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U68 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U69 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U70 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U71 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U72 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U73 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U74 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U75 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U76 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U77 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U78 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U79 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U80 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U81 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U82 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U83 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U84 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U85 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U86 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U87 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U88 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U89 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U90 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U91 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U92 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U93 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U94 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U95 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U96 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U97 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U98 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U99 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U100 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U101 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U102 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U103 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U104 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U105 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U106 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U107 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U108 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U109 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U110 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U111 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U112 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U113 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U114 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U115 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U116 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U117 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U118 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U119 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U120 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U121 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U122 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U123 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U124 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U125 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_25 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n197), .Z(result[9]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n194), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n193), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n193) );
  XOR2_X1 U134 ( .A(c[62]), .B(n192), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n191), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n190), .Z(result[60]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n188), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n187), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n186), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n185), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n184), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n183), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n182), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n181), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n180), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n179), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n178), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n177), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n176), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n175), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n174), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n173), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n172), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n171), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n170), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n169), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n168), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n167), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n166), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n165), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n164), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n163), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n162), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n161), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n160), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n159), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n158), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n157), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n156), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n155), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n154), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n153), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n152), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n151), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n150), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n149), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n148), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n147), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n146), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n145), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n144), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n143), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n142), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n141), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n140), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n139), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n138), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n137), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n136), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n135), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n134), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n196) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n195) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n194) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n192) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n191) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n190) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n188) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n187) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n186) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n185) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n184) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n183) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n182) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n181) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n180) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n179) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n177) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n167) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n176) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n175) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n174) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n173) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n172) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n171) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n170) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n169) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n168) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n166) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n156) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n165) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n164) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n163) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n162) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n161) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n160) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n159) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n158) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n157) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n155) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n145) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n154) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n153) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n152) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n151) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n150) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n149) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n148) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n147) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n146) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n144) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n134) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n143) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n142) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n141) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n140) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n139) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n138) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n137) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n136) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n135) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n197) );
  XOR2_X1 U2 ( .A(c[8]), .B(n196), .Z(result[8]) );
  INV_X1 U3 ( .A(c[5]), .ZN(n2) );
  INV_X1 U4 ( .A(a[4]), .ZN(n3) );
  INV_X1 U5 ( .A(a[5]), .ZN(n1) );
  XNOR2_X1 U6 ( .A(n1), .B(b[5]), .ZN(n189) );
  XNOR2_X1 U7 ( .A(n2), .B(n189), .ZN(result[5]) );
  XNOR2_X1 U8 ( .A(n3), .B(b[4]), .ZN(n178) );
  XOR2_X1 U9 ( .A(c[7]), .B(n195), .Z(result[7]) );
  AOI22_X1 U10 ( .A1(b[62]), .A2(a[62]), .B1(n192), .B2(c[62]), .ZN(n62) );
  INV_X1 U11 ( .A(n62), .ZN(carry[63]) );
  INV_X1 U12 ( .A(n12), .ZN(carry[18]) );
  AOI22_X1 U13 ( .A1(b[17]), .A2(a[17]), .B1(n142), .B2(c[17]), .ZN(n12) );
  INV_X1 U14 ( .A(n13), .ZN(carry[19]) );
  AOI22_X1 U15 ( .A1(b[18]), .A2(a[18]), .B1(n143), .B2(c[18]), .ZN(n13) );
  INV_X1 U16 ( .A(n6), .ZN(carry[12]) );
  AOI22_X1 U17 ( .A1(b[11]), .A2(a[11]), .B1(n136), .B2(c[11]), .ZN(n6) );
  INV_X1 U18 ( .A(n16), .ZN(carry[21]) );
  AOI22_X1 U19 ( .A1(b[20]), .A2(a[20]), .B1(n146), .B2(c[20]), .ZN(n16) );
  INV_X1 U20 ( .A(n15), .ZN(carry[20]) );
  AOI22_X1 U21 ( .A1(b[19]), .A2(a[19]), .B1(n144), .B2(c[19]), .ZN(n15) );
  INV_X1 U22 ( .A(n7), .ZN(carry[13]) );
  AOI22_X1 U23 ( .A1(b[12]), .A2(a[12]), .B1(n137), .B2(c[12]), .ZN(n7) );
  INV_X1 U24 ( .A(n11), .ZN(carry[17]) );
  AOI22_X1 U25 ( .A1(b[16]), .A2(a[16]), .B1(n141), .B2(c[16]), .ZN(n11) );
  INV_X1 U26 ( .A(n10), .ZN(carry[16]) );
  AOI22_X1 U27 ( .A1(b[15]), .A2(a[15]), .B1(n140), .B2(c[15]), .ZN(n10) );
  INV_X1 U28 ( .A(n8), .ZN(carry[14]) );
  AOI22_X1 U29 ( .A1(b[13]), .A2(a[13]), .B1(n138), .B2(c[13]), .ZN(n8) );
  INV_X1 U30 ( .A(n9), .ZN(carry[15]) );
  AOI22_X1 U31 ( .A1(b[14]), .A2(a[14]), .B1(n139), .B2(c[14]), .ZN(n9) );
  INV_X1 U32 ( .A(n17), .ZN(carry[22]) );
  AOI22_X1 U33 ( .A1(b[21]), .A2(a[21]), .B1(n147), .B2(c[21]), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(carry[23]) );
  AOI22_X1 U35 ( .A1(b[22]), .A2(a[22]), .B1(n148), .B2(c[22]), .ZN(n18) );
  INV_X1 U36 ( .A(n19), .ZN(carry[24]) );
  AOI22_X1 U37 ( .A1(b[23]), .A2(a[23]), .B1(n149), .B2(c[23]), .ZN(n19) );
  INV_X1 U38 ( .A(n20), .ZN(carry[25]) );
  AOI22_X1 U39 ( .A1(b[24]), .A2(a[24]), .B1(n150), .B2(c[24]), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(carry[26]) );
  AOI22_X1 U41 ( .A1(b[25]), .A2(a[25]), .B1(n151), .B2(c[25]), .ZN(n21) );
  INV_X1 U42 ( .A(n22), .ZN(carry[27]) );
  AOI22_X1 U43 ( .A1(b[26]), .A2(a[26]), .B1(n152), .B2(c[26]), .ZN(n22) );
  INV_X1 U44 ( .A(n23), .ZN(carry[28]) );
  AOI22_X1 U45 ( .A1(b[27]), .A2(a[27]), .B1(n153), .B2(c[27]), .ZN(n23) );
  INV_X1 U46 ( .A(n24), .ZN(carry[29]) );
  AOI22_X1 U47 ( .A1(b[28]), .A2(a[28]), .B1(n154), .B2(c[28]), .ZN(n24) );
  INV_X1 U48 ( .A(n26), .ZN(carry[30]) );
  AOI22_X1 U49 ( .A1(b[29]), .A2(a[29]), .B1(n155), .B2(c[29]), .ZN(n26) );
  INV_X1 U50 ( .A(n29), .ZN(carry[33]) );
  AOI22_X1 U51 ( .A1(b[32]), .A2(a[32]), .B1(n159), .B2(c[32]), .ZN(n29) );
  INV_X1 U52 ( .A(n30), .ZN(carry[34]) );
  AOI22_X1 U53 ( .A1(b[33]), .A2(a[33]), .B1(n160), .B2(c[33]), .ZN(n30) );
  INV_X1 U54 ( .A(n31), .ZN(carry[35]) );
  AOI22_X1 U55 ( .A1(b[34]), .A2(a[34]), .B1(n161), .B2(c[34]), .ZN(n31) );
  INV_X1 U56 ( .A(n32), .ZN(carry[36]) );
  AOI22_X1 U57 ( .A1(b[35]), .A2(a[35]), .B1(n162), .B2(c[35]), .ZN(n32) );
  INV_X1 U58 ( .A(n33), .ZN(carry[37]) );
  AOI22_X1 U59 ( .A1(b[36]), .A2(a[36]), .B1(n163), .B2(c[36]), .ZN(n33) );
  INV_X1 U60 ( .A(n34), .ZN(carry[38]) );
  AOI22_X1 U61 ( .A1(b[37]), .A2(a[37]), .B1(n164), .B2(c[37]), .ZN(n34) );
  INV_X1 U62 ( .A(n35), .ZN(carry[39]) );
  AOI22_X1 U63 ( .A1(b[38]), .A2(a[38]), .B1(n165), .B2(c[38]), .ZN(n35) );
  INV_X1 U64 ( .A(n37), .ZN(carry[40]) );
  AOI22_X1 U65 ( .A1(b[39]), .A2(a[39]), .B1(n166), .B2(c[39]), .ZN(n37) );
  INV_X1 U66 ( .A(n38), .ZN(carry[41]) );
  AOI22_X1 U67 ( .A1(b[40]), .A2(a[40]), .B1(n168), .B2(c[40]), .ZN(n38) );
  INV_X1 U68 ( .A(n39), .ZN(carry[42]) );
  AOI22_X1 U69 ( .A1(b[41]), .A2(a[41]), .B1(n169), .B2(c[41]), .ZN(n39) );
  INV_X1 U70 ( .A(n27), .ZN(carry[31]) );
  AOI22_X1 U71 ( .A1(b[30]), .A2(a[30]), .B1(n157), .B2(c[30]), .ZN(n27) );
  INV_X1 U72 ( .A(n28), .ZN(carry[32]) );
  AOI22_X1 U73 ( .A1(b[31]), .A2(a[31]), .B1(n158), .B2(c[31]), .ZN(n28) );
  INV_X1 U74 ( .A(n53), .ZN(carry[55]) );
  AOI22_X1 U75 ( .A1(b[54]), .A2(a[54]), .B1(n183), .B2(c[54]), .ZN(n53) );
  INV_X1 U76 ( .A(n40), .ZN(carry[43]) );
  AOI22_X1 U77 ( .A1(b[42]), .A2(a[42]), .B1(n170), .B2(c[42]), .ZN(n40) );
  INV_X1 U78 ( .A(n41), .ZN(carry[44]) );
  AOI22_X1 U79 ( .A1(b[43]), .A2(a[43]), .B1(n171), .B2(c[43]), .ZN(n41) );
  INV_X1 U80 ( .A(n42), .ZN(carry[45]) );
  AOI22_X1 U81 ( .A1(b[44]), .A2(a[44]), .B1(n172), .B2(c[44]), .ZN(n42) );
  INV_X1 U82 ( .A(n43), .ZN(carry[46]) );
  AOI22_X1 U83 ( .A1(b[45]), .A2(a[45]), .B1(n173), .B2(c[45]), .ZN(n43) );
  INV_X1 U84 ( .A(n44), .ZN(carry[47]) );
  AOI22_X1 U85 ( .A1(b[46]), .A2(a[46]), .B1(n174), .B2(c[46]), .ZN(n44) );
  INV_X1 U86 ( .A(n45), .ZN(carry[48]) );
  AOI22_X1 U87 ( .A1(b[47]), .A2(a[47]), .B1(n175), .B2(c[47]), .ZN(n45) );
  INV_X1 U88 ( .A(n46), .ZN(carry[49]) );
  AOI22_X1 U89 ( .A1(b[48]), .A2(a[48]), .B1(n176), .B2(c[48]), .ZN(n46) );
  INV_X1 U90 ( .A(n48), .ZN(carry[50]) );
  AOI22_X1 U91 ( .A1(b[49]), .A2(a[49]), .B1(n177), .B2(c[49]), .ZN(n48) );
  INV_X1 U92 ( .A(n49), .ZN(carry[51]) );
  AOI22_X1 U93 ( .A1(b[50]), .A2(a[50]), .B1(n179), .B2(c[50]), .ZN(n49) );
  INV_X1 U94 ( .A(n50), .ZN(carry[52]) );
  AOI22_X1 U95 ( .A1(b[51]), .A2(a[51]), .B1(n180), .B2(c[51]), .ZN(n50) );
  INV_X1 U96 ( .A(n51), .ZN(carry[53]) );
  AOI22_X1 U97 ( .A1(b[52]), .A2(a[52]), .B1(n181), .B2(c[52]), .ZN(n51) );
  INV_X1 U98 ( .A(n52), .ZN(carry[54]) );
  AOI22_X1 U99 ( .A1(b[53]), .A2(a[53]), .B1(n182), .B2(c[53]), .ZN(n52) );
  INV_X1 U100 ( .A(n57), .ZN(carry[59]) );
  AOI22_X1 U101 ( .A1(b[58]), .A2(a[58]), .B1(n187), .B2(c[58]), .ZN(n57) );
  INV_X1 U102 ( .A(n54), .ZN(carry[56]) );
  AOI22_X1 U103 ( .A1(b[55]), .A2(a[55]), .B1(n184), .B2(c[55]), .ZN(n54) );
  INV_X1 U104 ( .A(n55), .ZN(carry[57]) );
  AOI22_X1 U105 ( .A1(b[56]), .A2(a[56]), .B1(n185), .B2(c[56]), .ZN(n55) );
  INV_X1 U106 ( .A(n56), .ZN(carry[58]) );
  AOI22_X1 U107 ( .A1(b[57]), .A2(a[57]), .B1(n186), .B2(c[57]), .ZN(n56) );
  INV_X1 U108 ( .A(n59), .ZN(carry[60]) );
  AOI22_X1 U109 ( .A1(b[59]), .A2(a[59]), .B1(n188), .B2(c[59]), .ZN(n59) );
  INV_X1 U110 ( .A(n60), .ZN(carry[61]) );
  AOI22_X1 U111 ( .A1(b[60]), .A2(a[60]), .B1(n190), .B2(c[60]), .ZN(n60) );
  INV_X1 U112 ( .A(n61), .ZN(carry[62]) );
  AOI22_X1 U113 ( .A1(b[61]), .A2(a[61]), .B1(n191), .B2(c[61]), .ZN(n61) );
  INV_X1 U114 ( .A(n36), .ZN(carry[3]) );
  AOI22_X1 U115 ( .A1(b[2]), .A2(a[2]), .B1(n156), .B2(c[2]), .ZN(n36) );
  INV_X1 U116 ( .A(n47), .ZN(carry[4]) );
  AOI22_X1 U117 ( .A1(b[3]), .A2(a[3]), .B1(n167), .B2(c[3]), .ZN(n47) );
  INV_X1 U118 ( .A(n58), .ZN(carry[5]) );
  AOI22_X1 U119 ( .A1(b[4]), .A2(a[4]), .B1(n178), .B2(c[4]), .ZN(n58) );
  INV_X1 U120 ( .A(n63), .ZN(carry[6]) );
  AOI22_X1 U121 ( .A1(b[5]), .A2(a[5]), .B1(n189), .B2(c[5]), .ZN(n63) );
  INV_X1 U122 ( .A(n131), .ZN(carry[7]) );
  AOI22_X1 U123 ( .A1(b[6]), .A2(a[6]), .B1(n194), .B2(c[6]), .ZN(n131) );
  INV_X1 U124 ( .A(n132), .ZN(carry[8]) );
  AOI22_X1 U125 ( .A1(b[7]), .A2(a[7]), .B1(n195), .B2(c[7]), .ZN(n132) );
  INV_X1 U126 ( .A(n133), .ZN(carry[9]) );
  AOI22_X1 U127 ( .A1(b[8]), .A2(a[8]), .B1(n196), .B2(c[8]), .ZN(n133) );
  INV_X1 U129 ( .A(n4), .ZN(carry[10]) );
  AOI22_X1 U130 ( .A1(b[9]), .A2(a[9]), .B1(n197), .B2(c[9]), .ZN(n4) );
  INV_X1 U137 ( .A(n5), .ZN(carry[11]) );
  AOI22_X1 U196 ( .A1(b[10]), .A2(a[10]), .B1(n135), .B2(c[10]), .ZN(n5) );
  INV_X1 U201 ( .A(n25), .ZN(carry[2]) );
  AOI22_X1 U256 ( .A1(b[1]), .A2(a[1]), .B1(n145), .B2(c[1]), .ZN(n25) );
  INV_X1 U257 ( .A(n14), .ZN(carry[1]) );
  AOI22_X1 U258 ( .A1(b[0]), .A2(a[0]), .B1(n134), .B2(c[0]), .ZN(n14) );
endmodule


module BWAdder_26 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U3 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U4 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U5 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U6 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U7 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U8 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U9 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U10 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U11 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U12 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U13 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U14 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U15 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U16 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U17 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U18 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U19 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U20 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U21 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U22 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U23 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U24 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U25 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U26 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U27 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U28 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U29 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U30 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U31 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U32 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U33 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U34 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U35 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U36 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U37 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U38 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U39 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U40 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U41 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U42 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U43 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U44 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U45 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U46 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U47 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U48 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U49 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U50 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U51 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U52 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U53 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U54 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U55 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U56 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U57 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U58 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U59 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U60 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U61 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U62 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U63 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U64 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U65 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U66 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U67 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U68 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U69 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U70 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U71 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U72 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U73 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U74 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U75 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U76 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U77 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U78 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U79 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U80 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U81 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U82 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U83 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U84 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U85 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U86 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U87 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U88 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U89 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U90 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U91 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U92 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U93 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U94 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U95 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U96 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U97 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U98 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U99 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U100 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U101 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U102 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U103 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U104 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U105 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U106 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U107 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U108 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U109 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U110 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U111 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U112 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U113 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U114 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U115 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U116 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U117 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U118 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U119 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U120 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U121 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U122 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U123 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U124 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U125 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U126 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U127 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
endmodule


module BWAdder_27 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235;
  assign carry[0] = 1'b0;

  XOR2_X1 U132 ( .A(a[63]), .B(n231), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n231) );
  XOR2_X1 U134 ( .A(c[62]), .B(n230), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n229), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n228), .Z(result[60]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n226), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n225), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n224), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n223), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n222), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n221), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n220), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n219), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n218), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n217), .Z(result[50]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n215), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n214), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n213), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n212), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n211), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n210), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n209), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n208), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n207), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n206), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n205), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n204), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n203), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n202), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n201), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n200), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n199), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n198), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n197), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n196), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n195), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n194), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n193), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n192), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n191), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n190), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n189), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n188), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n187), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n186), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n185), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n184), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n183), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n182), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n181), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n180), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n179), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n178), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n177), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n176), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n175), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n174), .Z(result[11]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n172), .Z(result[0]) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n230) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n229) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n228) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n226) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n225) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n224) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n223) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n222) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n221) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n220) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n219) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n218) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n217) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n215) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n214) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n213) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n212) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n211) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n210) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n209) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n208) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n207) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n206) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n204) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n194) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n203) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n202) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n201) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n200) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n199) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n198) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n197) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n196) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n195) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n193) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n183) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n192) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n191) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n190) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n189) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n188) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n187) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n186) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n185) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n184) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n182) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n172) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n181) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n180) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n179) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n178) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n177) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n176) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n175) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n174) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n173) );
  INV_X1 U2 ( .A(n12), .ZN(n1) );
  INV_X1 U3 ( .A(c[10]), .ZN(n7) );
  INV_X1 U4 ( .A(c[4]), .ZN(n9) );
  INV_X1 U5 ( .A(c[5]), .ZN(n18) );
  INV_X1 U6 ( .A(c[7]), .ZN(n10) );
  INV_X1 U7 ( .A(c[8]), .ZN(n16) );
  INV_X1 U8 ( .A(c[9]), .ZN(n6) );
  INV_X1 U9 ( .A(b[3]), .ZN(n5) );
  INV_X1 U10 ( .A(b[4]), .ZN(n2) );
  INV_X1 U11 ( .A(b[5]), .ZN(n17) );
  INV_X1 U12 ( .A(b[6]), .ZN(n20) );
  INV_X1 U13 ( .A(b[7]), .ZN(n21) );
  INV_X1 U14 ( .A(b[8]), .ZN(n19) );
  XNOR2_X1 U15 ( .A(a[4]), .B(n2), .ZN(n216) );
  CLKBUF_X1 U16 ( .A(a[6]), .Z(n3) );
  CLKBUF_X1 U17 ( .A(n227), .Z(n4) );
  XNOR2_X1 U18 ( .A(a[3]), .B(n5), .ZN(n205) );
  XNOR2_X1 U19 ( .A(n235), .B(n6), .ZN(result[9]) );
  XNOR2_X1 U20 ( .A(n173), .B(n7), .ZN(result[10]) );
  CLKBUF_X1 U21 ( .A(a[8]), .Z(n8) );
  XNOR2_X1 U22 ( .A(n9), .B(n216), .ZN(result[4]) );
  XNOR2_X1 U23 ( .A(n233), .B(n10), .ZN(result[7]) );
  CLKBUF_X1 U24 ( .A(a[7]), .Z(n11) );
  NAND2_X1 U25 ( .A1(a[9]), .A2(n13), .ZN(n14) );
  NAND2_X1 U26 ( .A1(n12), .A2(b[9]), .ZN(n15) );
  NAND2_X1 U27 ( .A1(n15), .A2(n14), .ZN(n235) );
  INV_X1 U28 ( .A(a[9]), .ZN(n12) );
  INV_X1 U29 ( .A(b[9]), .ZN(n13) );
  XNOR2_X1 U30 ( .A(n234), .B(n16), .ZN(result[8]) );
  XNOR2_X1 U31 ( .A(a[5]), .B(n17), .ZN(n227) );
  XNOR2_X1 U32 ( .A(n227), .B(n18), .ZN(result[5]) );
  XNOR2_X1 U33 ( .A(a[8]), .B(n19), .ZN(n234) );
  XNOR2_X1 U34 ( .A(a[6]), .B(n20), .ZN(n232) );
  XNOR2_X1 U35 ( .A(a[7]), .B(n21), .ZN(n233) );
  INV_X1 U36 ( .A(n45), .ZN(carry[30]) );
  AOI22_X1 U37 ( .A1(b[29]), .A2(a[29]), .B1(n193), .B2(c[29]), .ZN(n45) );
  INV_X1 U38 ( .A(n41), .ZN(carry[27]) );
  AOI22_X1 U39 ( .A1(b[26]), .A2(a[26]), .B1(n190), .B2(c[26]), .ZN(n41) );
  INV_X1 U40 ( .A(n42), .ZN(carry[28]) );
  AOI22_X1 U41 ( .A1(b[27]), .A2(a[27]), .B1(n191), .B2(c[27]), .ZN(n42) );
  INV_X1 U42 ( .A(n43), .ZN(carry[29]) );
  AOI22_X1 U43 ( .A1(b[28]), .A2(a[28]), .B1(n192), .B2(c[28]), .ZN(n43) );
  INV_X1 U44 ( .A(n46), .ZN(carry[31]) );
  AOI22_X1 U45 ( .A1(b[30]), .A2(a[30]), .B1(n195), .B2(c[30]), .ZN(n46) );
  INV_X1 U46 ( .A(n47), .ZN(carry[32]) );
  AOI22_X1 U47 ( .A1(b[31]), .A2(a[31]), .B1(n196), .B2(c[31]), .ZN(n47) );
  INV_X1 U48 ( .A(n48), .ZN(carry[33]) );
  AOI22_X1 U49 ( .A1(b[32]), .A2(a[32]), .B1(n197), .B2(c[32]), .ZN(n48) );
  INV_X1 U50 ( .A(n49), .ZN(carry[34]) );
  AOI22_X1 U51 ( .A1(b[33]), .A2(a[33]), .B1(n198), .B2(c[33]), .ZN(n49) );
  INV_X1 U52 ( .A(n50), .ZN(carry[35]) );
  AOI22_X1 U53 ( .A1(b[34]), .A2(a[34]), .B1(n199), .B2(c[34]), .ZN(n50) );
  INV_X1 U54 ( .A(n51), .ZN(carry[36]) );
  AOI22_X1 U55 ( .A1(b[35]), .A2(a[35]), .B1(n200), .B2(c[35]), .ZN(n51) );
  INV_X1 U56 ( .A(n52), .ZN(carry[37]) );
  AOI22_X1 U57 ( .A1(b[36]), .A2(a[36]), .B1(n201), .B2(c[36]), .ZN(n52) );
  INV_X1 U58 ( .A(n53), .ZN(carry[38]) );
  AOI22_X1 U59 ( .A1(b[37]), .A2(a[37]), .B1(n202), .B2(c[37]), .ZN(n53) );
  INV_X1 U60 ( .A(n54), .ZN(carry[39]) );
  AOI22_X1 U61 ( .A1(b[38]), .A2(a[38]), .B1(n203), .B2(c[38]), .ZN(n54) );
  INV_X1 U62 ( .A(n56), .ZN(carry[40]) );
  AOI22_X1 U63 ( .A1(b[39]), .A2(a[39]), .B1(n204), .B2(c[39]), .ZN(n56) );
  INV_X1 U64 ( .A(n57), .ZN(carry[41]) );
  AOI22_X1 U65 ( .A1(b[40]), .A2(a[40]), .B1(n206), .B2(c[40]), .ZN(n57) );
  INV_X1 U66 ( .A(n58), .ZN(carry[42]) );
  AOI22_X1 U67 ( .A1(b[41]), .A2(a[41]), .B1(n207), .B2(c[41]), .ZN(n58) );
  INV_X1 U68 ( .A(n59), .ZN(carry[43]) );
  AOI22_X1 U69 ( .A1(b[42]), .A2(a[42]), .B1(n208), .B2(c[42]), .ZN(n59) );
  INV_X1 U70 ( .A(n60), .ZN(carry[44]) );
  AOI22_X1 U71 ( .A1(b[43]), .A2(a[43]), .B1(n209), .B2(c[43]), .ZN(n60) );
  INV_X1 U72 ( .A(n61), .ZN(carry[45]) );
  AOI22_X1 U73 ( .A1(b[44]), .A2(a[44]), .B1(n210), .B2(c[44]), .ZN(n61) );
  INV_X1 U74 ( .A(n62), .ZN(carry[46]) );
  AOI22_X1 U75 ( .A1(b[45]), .A2(a[45]), .B1(n211), .B2(c[45]), .ZN(n62) );
  INV_X1 U76 ( .A(n63), .ZN(carry[47]) );
  AOI22_X1 U77 ( .A1(b[46]), .A2(a[46]), .B1(n212), .B2(c[46]), .ZN(n63) );
  INV_X1 U78 ( .A(n150), .ZN(carry[48]) );
  AOI22_X1 U79 ( .A1(b[47]), .A2(a[47]), .B1(n213), .B2(c[47]), .ZN(n150) );
  INV_X1 U80 ( .A(n151), .ZN(carry[49]) );
  AOI22_X1 U81 ( .A1(b[48]), .A2(a[48]), .B1(n214), .B2(c[48]), .ZN(n151) );
  INV_X1 U82 ( .A(n153), .ZN(carry[50]) );
  AOI22_X1 U83 ( .A1(b[49]), .A2(a[49]), .B1(n215), .B2(c[49]), .ZN(n153) );
  INV_X1 U84 ( .A(n154), .ZN(carry[51]) );
  AOI22_X1 U85 ( .A1(b[50]), .A2(a[50]), .B1(n217), .B2(c[50]), .ZN(n154) );
  INV_X1 U86 ( .A(n155), .ZN(carry[52]) );
  AOI22_X1 U87 ( .A1(b[51]), .A2(a[51]), .B1(n218), .B2(c[51]), .ZN(n155) );
  INV_X1 U88 ( .A(n156), .ZN(carry[53]) );
  AOI22_X1 U89 ( .A1(b[52]), .A2(a[52]), .B1(n219), .B2(c[52]), .ZN(n156) );
  INV_X1 U90 ( .A(n157), .ZN(carry[54]) );
  AOI22_X1 U91 ( .A1(b[53]), .A2(a[53]), .B1(n220), .B2(c[53]), .ZN(n157) );
  INV_X1 U92 ( .A(n158), .ZN(carry[55]) );
  AOI22_X1 U93 ( .A1(b[54]), .A2(a[54]), .B1(n221), .B2(c[54]), .ZN(n158) );
  INV_X1 U94 ( .A(n159), .ZN(carry[56]) );
  AOI22_X1 U95 ( .A1(b[55]), .A2(a[55]), .B1(n222), .B2(c[55]), .ZN(n159) );
  INV_X1 U96 ( .A(n160), .ZN(carry[57]) );
  AOI22_X1 U97 ( .A1(b[56]), .A2(a[56]), .B1(n223), .B2(c[56]), .ZN(n160) );
  INV_X1 U98 ( .A(n161), .ZN(carry[58]) );
  AOI22_X1 U99 ( .A1(b[57]), .A2(a[57]), .B1(n224), .B2(c[57]), .ZN(n161) );
  INV_X1 U100 ( .A(n162), .ZN(carry[59]) );
  AOI22_X1 U101 ( .A1(b[58]), .A2(a[58]), .B1(n225), .B2(c[58]), .ZN(n162) );
  INV_X1 U102 ( .A(n164), .ZN(carry[60]) );
  AOI22_X1 U103 ( .A1(b[59]), .A2(a[59]), .B1(n226), .B2(c[59]), .ZN(n164) );
  INV_X1 U104 ( .A(n165), .ZN(carry[61]) );
  AOI22_X1 U105 ( .A1(b[60]), .A2(a[60]), .B1(n228), .B2(c[60]), .ZN(n165) );
  INV_X1 U106 ( .A(n166), .ZN(carry[62]) );
  AOI22_X1 U107 ( .A1(b[61]), .A2(a[61]), .B1(n229), .B2(c[61]), .ZN(n166) );
  INV_X1 U108 ( .A(n167), .ZN(carry[63]) );
  AOI22_X1 U109 ( .A1(b[62]), .A2(a[62]), .B1(n230), .B2(c[62]), .ZN(n167) );
  INV_X1 U110 ( .A(n24), .ZN(carry[11]) );
  INV_X1 U111 ( .A(n25), .ZN(carry[12]) );
  AOI22_X1 U112 ( .A1(b[11]), .A2(a[11]), .B1(n174), .B2(c[11]), .ZN(n25) );
  INV_X1 U113 ( .A(n26), .ZN(carry[13]) );
  AOI22_X1 U114 ( .A1(b[12]), .A2(a[12]), .B1(n175), .B2(c[12]), .ZN(n26) );
  INV_X1 U115 ( .A(n27), .ZN(carry[14]) );
  AOI22_X1 U116 ( .A1(b[13]), .A2(a[13]), .B1(n176), .B2(c[13]), .ZN(n27) );
  INV_X1 U117 ( .A(c[6]), .ZN(n22) );
  INV_X1 U118 ( .A(n23), .ZN(carry[10]) );
  INV_X1 U119 ( .A(n36), .ZN(carry[22]) );
  AOI22_X1 U120 ( .A1(b[21]), .A2(a[21]), .B1(n185), .B2(c[21]), .ZN(n36) );
  INV_X1 U121 ( .A(n35), .ZN(carry[21]) );
  AOI22_X1 U122 ( .A1(b[20]), .A2(a[20]), .B1(n184), .B2(c[20]), .ZN(n35) );
  INV_X1 U123 ( .A(n34), .ZN(carry[20]) );
  AOI22_X1 U124 ( .A1(b[19]), .A2(a[19]), .B1(n182), .B2(c[19]), .ZN(n34) );
  INV_X1 U125 ( .A(n32), .ZN(carry[19]) );
  AOI22_X1 U126 ( .A1(b[18]), .A2(a[18]), .B1(n181), .B2(c[18]), .ZN(n32) );
  INV_X1 U127 ( .A(n37), .ZN(carry[23]) );
  AOI22_X1 U128 ( .A1(b[22]), .A2(a[22]), .B1(n186), .B2(c[22]), .ZN(n37) );
  INV_X1 U129 ( .A(n38), .ZN(carry[24]) );
  AOI22_X1 U130 ( .A1(b[23]), .A2(a[23]), .B1(n187), .B2(c[23]), .ZN(n38) );
  INV_X1 U131 ( .A(n39), .ZN(carry[25]) );
  AOI22_X1 U137 ( .A1(b[24]), .A2(a[24]), .B1(n188), .B2(c[24]), .ZN(n39) );
  INV_X1 U148 ( .A(n40), .ZN(carry[26]) );
  AOI22_X1 U191 ( .A1(b[25]), .A2(a[25]), .B1(n189), .B2(c[25]), .ZN(n40) );
  INV_X1 U193 ( .A(n30), .ZN(carry[17]) );
  AOI22_X1 U194 ( .A1(b[16]), .A2(a[16]), .B1(n179), .B2(c[16]), .ZN(n30) );
  INV_X1 U195 ( .A(n29), .ZN(carry[16]) );
  AOI22_X1 U196 ( .A1(b[15]), .A2(a[15]), .B1(n178), .B2(c[15]), .ZN(n29) );
  INV_X1 U201 ( .A(n31), .ZN(carry[18]) );
  AOI22_X1 U212 ( .A1(b[17]), .A2(a[17]), .B1(n180), .B2(c[17]), .ZN(n31) );
  INV_X1 U255 ( .A(n28), .ZN(carry[15]) );
  AOI22_X1 U256 ( .A1(b[14]), .A2(a[14]), .B1(n177), .B2(c[14]), .ZN(n28) );
  INV_X1 U257 ( .A(n169), .ZN(carry[7]) );
  INV_X1 U258 ( .A(n152), .ZN(carry[4]) );
  INV_X1 U259 ( .A(n163), .ZN(carry[5]) );
  INV_X1 U260 ( .A(n168), .ZN(carry[6]) );
  INV_X1 U261 ( .A(n170), .ZN(carry[8]) );
  INV_X1 U262 ( .A(n171), .ZN(carry[9]) );
  INV_X1 U263 ( .A(n33), .ZN(carry[1]) );
  AOI22_X1 U264 ( .A1(b[0]), .A2(a[0]), .B1(n172), .B2(c[0]), .ZN(n33) );
  INV_X1 U265 ( .A(n44), .ZN(carry[2]) );
  AOI22_X1 U266 ( .A1(b[1]), .A2(a[1]), .B1(n183), .B2(c[1]), .ZN(n44) );
  INV_X1 U267 ( .A(n55), .ZN(carry[3]) );
  AOI22_X1 U268 ( .A1(b[2]), .A2(a[2]), .B1(n194), .B2(c[2]), .ZN(n55) );
  AOI22_X1 U269 ( .A1(b[7]), .A2(n11), .B1(n233), .B2(c[7]), .ZN(n170) );
  AOI22_X1 U270 ( .A1(b[3]), .A2(a[3]), .B1(n205), .B2(c[3]), .ZN(n152) );
  XNOR2_X1 U271 ( .A(n232), .B(n22), .ZN(result[6]) );
  AOI22_X1 U272 ( .A1(b[4]), .A2(a[4]), .B1(n216), .B2(c[4]), .ZN(n163) );
  AOI22_X1 U273 ( .A1(b[10]), .A2(a[10]), .B1(n173), .B2(c[10]), .ZN(n24) );
  AOI22_X1 U274 ( .A1(b[9]), .A2(n1), .B1(n235), .B2(c[9]), .ZN(n23) );
  AOI22_X1 U275 ( .A1(b[8]), .A2(n8), .B1(n234), .B2(c[8]), .ZN(n171) );
  AOI22_X1 U276 ( .A1(b[5]), .A2(a[5]), .B1(n4), .B2(c[5]), .ZN(n168) );
  AOI22_X1 U277 ( .A1(b[6]), .A2(n3), .B1(n232), .B2(c[6]), .ZN(n169) );
endmodule


module BWAdder_28 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U3 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U4 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U5 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U6 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U7 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U8 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U9 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U10 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U11 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U12 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U13 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U14 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U15 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U16 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U17 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U18 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U19 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U20 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U21 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U22 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U23 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U24 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U25 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U26 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U27 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U28 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U29 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U30 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U31 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U32 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U33 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U34 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U35 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U36 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U37 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U38 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U39 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U40 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U41 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U42 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U43 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U44 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U45 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U46 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U47 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U48 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U49 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U50 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U51 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U52 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U53 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U54 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U55 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U56 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U57 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U58 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U59 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U60 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U61 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U62 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U63 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U64 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U65 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U66 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U67 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U68 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U69 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U70 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U71 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U72 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U73 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U74 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U75 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U76 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U77 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U78 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U79 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U80 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U81 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U82 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U83 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U84 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U85 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U86 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U87 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U88 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U89 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U90 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U91 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U92 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U93 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U94 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U95 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U96 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U97 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U98 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U99 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U100 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U101 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U102 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U103 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U104 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U105 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U106 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U107 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U108 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U109 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U110 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U111 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U112 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U113 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U114 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U115 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U116 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U117 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U118 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U119 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U120 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U121 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U122 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U123 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U124 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U125 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_29 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U3 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U4 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U5 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U6 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U7 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U8 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U9 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U10 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U11 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U12 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U13 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U14 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U15 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U16 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U17 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U18 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U19 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U20 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U21 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U22 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U23 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U24 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U25 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U26 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U27 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U28 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U29 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U30 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U31 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U32 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U33 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U34 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U35 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U36 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U37 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U38 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U39 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U40 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U41 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U42 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U43 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U44 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U45 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U46 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U47 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U48 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U49 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U50 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U51 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U52 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U53 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U54 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U55 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U56 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U57 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U58 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U59 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U60 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U61 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U62 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U63 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U64 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U65 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U66 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U67 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U68 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U69 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U70 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U71 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U72 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U73 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U74 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U75 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U76 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U77 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U78 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U79 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U80 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U81 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U82 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U83 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U84 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U85 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U86 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U87 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U88 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U89 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U90 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U91 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U92 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U93 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U94 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U95 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U96 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U97 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U98 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U99 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U100 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U101 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U102 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U103 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U104 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U105 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U106 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U107 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U108 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U109 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U110 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U111 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U112 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U113 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U114 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U115 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U116 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U117 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U118 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U119 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U120 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U121 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U122 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U123 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U124 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U125 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_30 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U3 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U4 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U5 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U6 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U7 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U8 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U9 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U10 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U11 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U12 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U13 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U14 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U15 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U16 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U17 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U18 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U19 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U20 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U21 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U22 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U23 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U24 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U25 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U26 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U27 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U28 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U29 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U30 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U31 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U32 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U33 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U34 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U35 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U36 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U37 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U38 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U39 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U40 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U41 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U42 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U43 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U44 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U45 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U46 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U47 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U48 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U49 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U50 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U51 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U52 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U53 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U54 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U55 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U56 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U57 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U58 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U59 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U60 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U61 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U62 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U63 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U64 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U65 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U66 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U67 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U68 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U69 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U70 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U71 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U72 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U73 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U74 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U75 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U76 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U77 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U78 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U79 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U80 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U81 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U82 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U83 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U84 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U85 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U86 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U87 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U88 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U89 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U90 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U91 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U92 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U93 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U94 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U95 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U96 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U97 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U98 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U99 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U100 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U101 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U102 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U103 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U104 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U105 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U106 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U107 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U108 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U109 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U110 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U111 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U112 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U113 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U114 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U115 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U116 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U117 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U118 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U119 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U120 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U121 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U122 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U123 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U124 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U125 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_31 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U3 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U4 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U5 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U6 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U7 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U8 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U9 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U10 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U11 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U12 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U13 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U14 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U15 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U16 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U17 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U18 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U19 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U20 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U21 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U22 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U23 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U24 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U25 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U26 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U27 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U28 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U29 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U30 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U31 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U32 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U33 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U34 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U35 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U36 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U37 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U38 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U39 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U40 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U41 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U42 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U43 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U44 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U45 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U46 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U47 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U48 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U49 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U50 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U51 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U52 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U53 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U54 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U55 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U56 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U57 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U58 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U59 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U60 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U61 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U62 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U63 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U64 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U65 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U66 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U67 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U68 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U69 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U70 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U71 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U72 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U73 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U74 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U75 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U76 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U77 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U78 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U79 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U80 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U81 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U82 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U83 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U84 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U85 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U86 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U87 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U88 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U89 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U90 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U91 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U92 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U93 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U94 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U95 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U96 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U97 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U98 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U99 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U100 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U101 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U102 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U103 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U104 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U105 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U106 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U107 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U108 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U109 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U110 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U111 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U112 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U113 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U114 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U115 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U116 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U117 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U118 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U119 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U120 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U121 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U122 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U123 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U124 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U125 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_32 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U3 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U4 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U5 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U6 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U7 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U8 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U9 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U10 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U11 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U12 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U13 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U14 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U15 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U16 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U17 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U18 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U19 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U20 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U21 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U22 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U23 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U24 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U25 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U26 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U27 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U28 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U29 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U30 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U31 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U32 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U33 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U34 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U35 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U36 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U37 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U38 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U39 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U40 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U41 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U42 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U43 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U44 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U45 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U46 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U47 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U48 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U49 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U50 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U51 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U52 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U53 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U54 ( .A(n59), .ZN(carry[63]) );
  INV_X1 U55 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U56 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U57 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U58 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U59 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U60 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U61 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U62 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U63 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U64 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U65 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U66 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U67 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U68 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U69 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U70 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U71 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U72 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  AOI22_X1 U73 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U74 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U75 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U76 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U77 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U78 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U79 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U80 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U81 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U82 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U83 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U84 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U85 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U86 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U87 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U88 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U89 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U90 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U91 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U92 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U93 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U94 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U95 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U96 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U97 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U98 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U99 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U100 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U101 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U102 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U103 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U104 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U105 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U106 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U107 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U108 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U109 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U110 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U111 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U112 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U113 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U114 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U115 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U116 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U117 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U118 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U119 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U120 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U121 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U122 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U123 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U124 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U125 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_33 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U3 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U4 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U5 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U6 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U7 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U8 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U9 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U10 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U11 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U12 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U13 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U14 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U15 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U16 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U17 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U18 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U19 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U20 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U21 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U22 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U23 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U24 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U25 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U26 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U27 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U28 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U29 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U30 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U31 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U32 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U33 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U34 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U35 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U36 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U37 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U38 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U39 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U40 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U41 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U42 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U43 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U44 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U45 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U46 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U47 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U48 ( .A(n59), .ZN(carry[63]) );
  INV_X1 U49 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U50 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U51 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U52 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U53 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U54 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U55 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U56 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U57 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U58 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U59 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U60 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U61 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U62 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U63 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U64 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U65 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U66 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U67 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U68 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U69 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U70 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U71 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U72 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U73 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U74 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U75 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U76 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U77 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U78 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U79 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U80 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U81 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U82 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U83 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U84 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U85 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U86 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U87 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U88 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U89 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U90 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  AOI22_X1 U91 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U92 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U93 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U94 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U95 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U96 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U97 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U98 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U99 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U100 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U101 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U102 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U103 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U104 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U105 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U106 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U107 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U108 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U109 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U110 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U111 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U112 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U113 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U114 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U115 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U116 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U117 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U118 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U119 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U120 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U121 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U122 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U123 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U124 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U125 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U126 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U127 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
endmodule


module BWAdder_34 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n193), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n192), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n191), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n190), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n189), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n189) );
  XOR2_X1 U134 ( .A(c[62]), .B(n188), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n187), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n186), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n185), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n184), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n183), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n182), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n181), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n180), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n179), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n178), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n177), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n176), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n175), .Z(result[50]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n173), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n172), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n171), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n170), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n169), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n168), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n167), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n166), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n165), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n164), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n163), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n162), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n161), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n160), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n159), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n158), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n157), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n156), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n155), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n154), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n153), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n152), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n151), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n150), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n149), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n148), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n147), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n146), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n145), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n144), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n143), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n142), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n141), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n140), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n139), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n138), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n137), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n136), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n135), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n134), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n133), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n132), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n131), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n130), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n192) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n191) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n190) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n185) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n188) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n187) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n186) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n184) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n174) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n183) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n182) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n181) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n180) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n179) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n178) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n177) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n176) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n175) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n173) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n163) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n172) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n171) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n170) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n169) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n168) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n167) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n166) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n165) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n164) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n162) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n152) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n161) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n160) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n159) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n158) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n157) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n156) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n155) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n154) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n153) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n151) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n141) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n150) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n149) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n148) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n147) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n146) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n145) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n144) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n143) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n142) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n140) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n130) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n139) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n138) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n137) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n136) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n135) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n134) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n133) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n132) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n131) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n193) );
  INV_X1 U2 ( .A(c[4]), .ZN(n1) );
  XNOR2_X1 U3 ( .A(n1), .B(n174), .ZN(result[4]) );
  INV_X1 U4 ( .A(n15), .ZN(carry[22]) );
  AOI22_X1 U5 ( .A1(b[21]), .A2(a[21]), .B1(n143), .B2(c[21]), .ZN(n15) );
  INV_X1 U6 ( .A(n16), .ZN(carry[23]) );
  AOI22_X1 U7 ( .A1(b[22]), .A2(a[22]), .B1(n144), .B2(c[22]), .ZN(n16) );
  INV_X1 U8 ( .A(n17), .ZN(carry[24]) );
  AOI22_X1 U9 ( .A1(b[23]), .A2(a[23]), .B1(n145), .B2(c[23]), .ZN(n17) );
  INV_X1 U10 ( .A(n18), .ZN(carry[25]) );
  AOI22_X1 U11 ( .A1(b[24]), .A2(a[24]), .B1(n146), .B2(c[24]), .ZN(n18) );
  INV_X1 U12 ( .A(n19), .ZN(carry[26]) );
  AOI22_X1 U13 ( .A1(b[25]), .A2(a[25]), .B1(n147), .B2(c[25]), .ZN(n19) );
  INV_X1 U14 ( .A(n20), .ZN(carry[27]) );
  AOI22_X1 U15 ( .A1(b[26]), .A2(a[26]), .B1(n148), .B2(c[26]), .ZN(n20) );
  INV_X1 U16 ( .A(n21), .ZN(carry[28]) );
  AOI22_X1 U17 ( .A1(b[27]), .A2(a[27]), .B1(n149), .B2(c[27]), .ZN(n21) );
  INV_X1 U18 ( .A(n22), .ZN(carry[29]) );
  AOI22_X1 U19 ( .A1(b[28]), .A2(a[28]), .B1(n150), .B2(c[28]), .ZN(n22) );
  INV_X1 U20 ( .A(n24), .ZN(carry[30]) );
  AOI22_X1 U21 ( .A1(b[29]), .A2(a[29]), .B1(n151), .B2(c[29]), .ZN(n24) );
  INV_X1 U22 ( .A(n13), .ZN(carry[20]) );
  AOI22_X1 U23 ( .A1(b[19]), .A2(a[19]), .B1(n140), .B2(c[19]), .ZN(n13) );
  INV_X1 U24 ( .A(n11), .ZN(carry[19]) );
  AOI22_X1 U25 ( .A1(b[18]), .A2(a[18]), .B1(n139), .B2(c[18]), .ZN(n11) );
  INV_X1 U26 ( .A(n10), .ZN(carry[18]) );
  AOI22_X1 U27 ( .A1(b[17]), .A2(a[17]), .B1(n138), .B2(c[17]), .ZN(n10) );
  INV_X1 U28 ( .A(n9), .ZN(carry[17]) );
  AOI22_X1 U29 ( .A1(b[16]), .A2(a[16]), .B1(n137), .B2(c[16]), .ZN(n9) );
  INV_X1 U30 ( .A(n14), .ZN(carry[21]) );
  AOI22_X1 U31 ( .A1(b[20]), .A2(a[20]), .B1(n142), .B2(c[20]), .ZN(n14) );
  INV_X1 U32 ( .A(n4), .ZN(carry[12]) );
  AOI22_X1 U33 ( .A1(b[11]), .A2(a[11]), .B1(n132), .B2(c[11]), .ZN(n4) );
  INV_X1 U34 ( .A(n5), .ZN(carry[13]) );
  AOI22_X1 U35 ( .A1(b[12]), .A2(a[12]), .B1(n133), .B2(c[12]), .ZN(n5) );
  INV_X1 U36 ( .A(n6), .ZN(carry[14]) );
  AOI22_X1 U37 ( .A1(b[13]), .A2(a[13]), .B1(n134), .B2(c[13]), .ZN(n6) );
  INV_X1 U38 ( .A(n7), .ZN(carry[15]) );
  AOI22_X1 U39 ( .A1(b[14]), .A2(a[14]), .B1(n135), .B2(c[14]), .ZN(n7) );
  INV_X1 U40 ( .A(n8), .ZN(carry[16]) );
  AOI22_X1 U41 ( .A1(b[15]), .A2(a[15]), .B1(n136), .B2(c[15]), .ZN(n8) );
  INV_X1 U42 ( .A(n25), .ZN(carry[31]) );
  AOI22_X1 U43 ( .A1(b[30]), .A2(a[30]), .B1(n153), .B2(c[30]), .ZN(n25) );
  INV_X1 U44 ( .A(n2), .ZN(carry[10]) );
  AOI22_X1 U45 ( .A1(b[9]), .A2(a[9]), .B1(n193), .B2(c[9]), .ZN(n2) );
  INV_X1 U46 ( .A(n3), .ZN(carry[11]) );
  AOI22_X1 U47 ( .A1(b[10]), .A2(a[10]), .B1(n131), .B2(c[10]), .ZN(n3) );
  INV_X1 U48 ( .A(n27), .ZN(carry[33]) );
  AOI22_X1 U49 ( .A1(b[32]), .A2(a[32]), .B1(n155), .B2(c[32]), .ZN(n27) );
  INV_X1 U50 ( .A(n28), .ZN(carry[34]) );
  AOI22_X1 U51 ( .A1(b[33]), .A2(a[33]), .B1(n156), .B2(c[33]), .ZN(n28) );
  INV_X1 U52 ( .A(n29), .ZN(carry[35]) );
  AOI22_X1 U53 ( .A1(b[34]), .A2(a[34]), .B1(n157), .B2(c[34]), .ZN(n29) );
  INV_X1 U54 ( .A(n30), .ZN(carry[36]) );
  AOI22_X1 U55 ( .A1(b[35]), .A2(a[35]), .B1(n158), .B2(c[35]), .ZN(n30) );
  INV_X1 U56 ( .A(n31), .ZN(carry[37]) );
  AOI22_X1 U57 ( .A1(b[36]), .A2(a[36]), .B1(n159), .B2(c[36]), .ZN(n31) );
  INV_X1 U58 ( .A(n32), .ZN(carry[38]) );
  AOI22_X1 U59 ( .A1(b[37]), .A2(a[37]), .B1(n160), .B2(c[37]), .ZN(n32) );
  INV_X1 U60 ( .A(n33), .ZN(carry[39]) );
  AOI22_X1 U61 ( .A1(b[38]), .A2(a[38]), .B1(n161), .B2(c[38]), .ZN(n33) );
  INV_X1 U62 ( .A(n35), .ZN(carry[40]) );
  AOI22_X1 U63 ( .A1(b[39]), .A2(a[39]), .B1(n162), .B2(c[39]), .ZN(n35) );
  INV_X1 U64 ( .A(n36), .ZN(carry[41]) );
  AOI22_X1 U65 ( .A1(b[40]), .A2(a[40]), .B1(n164), .B2(c[40]), .ZN(n36) );
  INV_X1 U66 ( .A(n37), .ZN(carry[42]) );
  AOI22_X1 U67 ( .A1(b[41]), .A2(a[41]), .B1(n165), .B2(c[41]), .ZN(n37) );
  INV_X1 U68 ( .A(n26), .ZN(carry[32]) );
  AOI22_X1 U69 ( .A1(b[31]), .A2(a[31]), .B1(n154), .B2(c[31]), .ZN(n26) );
  INV_X1 U70 ( .A(n43), .ZN(carry[48]) );
  AOI22_X1 U71 ( .A1(b[47]), .A2(a[47]), .B1(n171), .B2(c[47]), .ZN(n43) );
  INV_X1 U72 ( .A(n46), .ZN(carry[50]) );
  AOI22_X1 U73 ( .A1(b[49]), .A2(a[49]), .B1(n173), .B2(c[49]), .ZN(n46) );
  INV_X1 U74 ( .A(n48), .ZN(carry[52]) );
  AOI22_X1 U75 ( .A1(b[51]), .A2(a[51]), .B1(n176), .B2(c[51]), .ZN(n48) );
  INV_X1 U76 ( .A(n51), .ZN(carry[55]) );
  AOI22_X1 U77 ( .A1(b[54]), .A2(a[54]), .B1(n179), .B2(c[54]), .ZN(n51) );
  INV_X1 U78 ( .A(n38), .ZN(carry[43]) );
  AOI22_X1 U79 ( .A1(b[42]), .A2(a[42]), .B1(n166), .B2(c[42]), .ZN(n38) );
  INV_X1 U80 ( .A(n39), .ZN(carry[44]) );
  AOI22_X1 U81 ( .A1(b[43]), .A2(a[43]), .B1(n167), .B2(c[43]), .ZN(n39) );
  INV_X1 U82 ( .A(n40), .ZN(carry[45]) );
  AOI22_X1 U83 ( .A1(b[44]), .A2(a[44]), .B1(n168), .B2(c[44]), .ZN(n40) );
  INV_X1 U84 ( .A(n41), .ZN(carry[46]) );
  AOI22_X1 U85 ( .A1(b[45]), .A2(a[45]), .B1(n169), .B2(c[45]), .ZN(n41) );
  INV_X1 U86 ( .A(n42), .ZN(carry[47]) );
  AOI22_X1 U87 ( .A1(b[46]), .A2(a[46]), .B1(n170), .B2(c[46]), .ZN(n42) );
  INV_X1 U88 ( .A(n44), .ZN(carry[49]) );
  AOI22_X1 U89 ( .A1(b[48]), .A2(a[48]), .B1(n172), .B2(c[48]), .ZN(n44) );
  INV_X1 U90 ( .A(n47), .ZN(carry[51]) );
  AOI22_X1 U91 ( .A1(b[50]), .A2(a[50]), .B1(n175), .B2(c[50]), .ZN(n47) );
  INV_X1 U92 ( .A(n49), .ZN(carry[53]) );
  AOI22_X1 U93 ( .A1(b[52]), .A2(a[52]), .B1(n177), .B2(c[52]), .ZN(n49) );
  INV_X1 U94 ( .A(n50), .ZN(carry[54]) );
  AOI22_X1 U95 ( .A1(b[53]), .A2(a[53]), .B1(n178), .B2(c[53]), .ZN(n50) );
  INV_X1 U96 ( .A(n52), .ZN(carry[56]) );
  AOI22_X1 U97 ( .A1(b[55]), .A2(a[55]), .B1(n180), .B2(c[55]), .ZN(n52) );
  INV_X1 U98 ( .A(n54), .ZN(carry[58]) );
  AOI22_X1 U99 ( .A1(b[57]), .A2(a[57]), .B1(n182), .B2(c[57]), .ZN(n54) );
  INV_X1 U100 ( .A(n55), .ZN(carry[59]) );
  AOI22_X1 U101 ( .A1(b[58]), .A2(a[58]), .B1(n183), .B2(c[58]), .ZN(n55) );
  INV_X1 U102 ( .A(n57), .ZN(carry[60]) );
  AOI22_X1 U103 ( .A1(b[59]), .A2(a[59]), .B1(n184), .B2(c[59]), .ZN(n57) );
  INV_X1 U104 ( .A(n53), .ZN(carry[57]) );
  AOI22_X1 U105 ( .A1(b[56]), .A2(a[56]), .B1(n181), .B2(c[56]), .ZN(n53) );
  INV_X1 U106 ( .A(n58), .ZN(carry[61]) );
  AOI22_X1 U107 ( .A1(b[60]), .A2(a[60]), .B1(n186), .B2(c[60]), .ZN(n58) );
  INV_X1 U108 ( .A(n59), .ZN(carry[62]) );
  AOI22_X1 U109 ( .A1(b[61]), .A2(a[61]), .B1(n187), .B2(c[61]), .ZN(n59) );
  INV_X1 U110 ( .A(n60), .ZN(carry[63]) );
  AOI22_X1 U111 ( .A1(b[62]), .A2(a[62]), .B1(n188), .B2(c[62]), .ZN(n60) );
  INV_X1 U112 ( .A(n61), .ZN(carry[6]) );
  AOI22_X1 U113 ( .A1(b[5]), .A2(a[5]), .B1(n185), .B2(c[5]), .ZN(n61) );
  INV_X1 U114 ( .A(n129), .ZN(carry[9]) );
  AOI22_X1 U115 ( .A1(b[8]), .A2(a[8]), .B1(n192), .B2(c[8]), .ZN(n129) );
  INV_X1 U116 ( .A(n63), .ZN(carry[8]) );
  AOI22_X1 U117 ( .A1(b[7]), .A2(a[7]), .B1(n191), .B2(c[7]), .ZN(n63) );
  INV_X1 U118 ( .A(n62), .ZN(carry[7]) );
  AOI22_X1 U119 ( .A1(b[6]), .A2(a[6]), .B1(n190), .B2(c[6]), .ZN(n62) );
  INV_X1 U120 ( .A(n34), .ZN(carry[3]) );
  AOI22_X1 U121 ( .A1(b[2]), .A2(a[2]), .B1(n152), .B2(c[2]), .ZN(n34) );
  INV_X1 U122 ( .A(n45), .ZN(carry[4]) );
  AOI22_X1 U123 ( .A1(b[3]), .A2(a[3]), .B1(n163), .B2(c[3]), .ZN(n45) );
  INV_X1 U124 ( .A(n56), .ZN(carry[5]) );
  AOI22_X1 U125 ( .A1(b[4]), .A2(a[4]), .B1(n174), .B2(c[4]), .ZN(n56) );
  INV_X1 U126 ( .A(n23), .ZN(carry[2]) );
  AOI22_X1 U127 ( .A1(b[1]), .A2(a[1]), .B1(n141), .B2(c[1]), .ZN(n23) );
  INV_X1 U148 ( .A(n12), .ZN(carry[1]) );
  AOI22_X1 U256 ( .A1(b[0]), .A2(a[0]), .B1(n130), .B2(c[0]), .ZN(n12) );
endmodule


module BWAdder_35 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U3 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U4 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U5 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U6 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U7 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U8 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U9 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U10 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U11 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U12 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U13 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U14 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U15 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U16 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U17 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U18 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U19 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U20 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U21 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U22 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U23 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U24 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U25 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U26 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U27 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U28 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U29 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U30 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U31 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U32 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U33 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U34 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U35 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U36 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U37 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U38 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U39 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U40 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U41 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U42 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U43 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U44 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U45 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U46 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U47 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U48 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U49 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U50 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U51 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U52 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U53 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U54 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U55 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U56 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U57 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U58 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U59 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U60 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U61 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U62 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U63 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U64 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U65 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U66 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U67 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U68 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U69 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U70 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U71 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U72 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U73 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U74 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U75 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U76 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U77 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U78 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U79 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U80 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U81 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U82 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U83 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U84 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U85 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U86 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U87 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U88 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U89 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U90 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U91 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U92 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U93 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U94 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U95 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U96 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U97 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U98 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U99 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U100 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U101 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U102 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U103 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U104 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U105 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U106 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U107 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U108 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U109 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U110 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U111 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U112 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U113 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U114 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U115 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U116 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U117 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U118 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U119 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U120 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U121 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U122 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U123 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U124 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U125 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U126 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U127 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
endmodule


module BWAdder_36 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U3 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U4 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U5 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U6 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U7 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U8 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U9 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U10 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U11 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U12 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U13 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U14 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U15 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U16 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U17 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U18 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U19 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  AOI22_X1 U20 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U21 ( .A(n59), .ZN(carry[63]) );
  INV_X1 U22 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U23 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U24 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U25 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U26 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U27 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U28 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U29 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U30 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U31 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U32 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U33 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U34 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U35 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U36 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U37 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U38 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U39 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U40 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U41 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U42 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U43 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U44 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U45 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U46 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U47 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U48 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U49 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U50 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U51 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U52 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U53 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U54 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U55 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U56 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U57 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U58 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U59 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U60 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U61 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U62 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U63 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U64 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U65 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U66 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U67 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U68 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U69 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U70 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U71 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U72 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U73 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U74 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U75 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U76 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U77 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U78 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U79 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U80 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U81 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U82 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U83 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U84 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U85 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U86 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U87 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U88 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U89 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U90 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U91 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U92 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U93 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U94 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U95 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U96 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U97 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U98 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U99 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U100 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U101 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U102 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U103 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U104 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U105 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U106 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U107 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U108 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U109 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U110 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U111 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U112 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U113 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U114 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U115 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U116 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U117 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U118 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U119 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U120 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U121 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U122 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U123 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U124 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U125 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U126 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U127 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
endmodule


module BWAdder_37 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U3 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U4 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U5 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U6 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U7 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U8 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U9 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U10 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U11 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U12 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U13 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U14 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U15 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U16 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U17 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U18 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U19 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U20 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U21 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U22 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U23 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U24 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U25 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U26 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U27 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U28 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U29 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U30 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U31 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U32 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U33 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U34 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U35 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U36 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U37 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U38 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U39 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U40 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U41 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U42 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U43 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U44 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U45 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U46 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U47 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U48 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U49 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U50 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U51 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U52 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U53 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U54 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U55 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U56 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U57 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U58 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U59 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U60 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U61 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U62 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U63 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U64 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U65 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U66 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U67 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U68 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U69 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U70 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U72 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U73 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U74 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U75 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U76 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U77 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U78 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U79 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U80 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U81 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U82 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U83 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U84 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U85 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U86 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U87 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U88 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U89 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U90 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U91 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U92 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U93 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U94 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U95 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U96 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U97 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U98 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U99 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U100 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U101 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U102 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U103 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U104 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U105 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U106 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U107 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U108 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U109 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U110 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U111 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U112 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U113 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U114 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U115 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U116 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U117 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U118 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U119 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U120 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U121 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U122 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U123 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U124 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U125 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U126 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U127 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
endmodule


module BWAdder_38 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U3 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U4 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U5 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U6 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U7 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U8 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U9 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U10 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U11 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U12 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U13 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U14 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U15 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U16 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U17 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U18 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U19 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U20 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U21 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U22 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U23 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U24 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U25 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U26 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U27 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U28 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U29 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U30 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U31 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U32 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U33 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U34 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U35 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U36 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U37 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U38 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U39 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U40 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U41 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U42 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U43 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U44 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U45 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U46 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U47 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U48 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U49 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U50 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U51 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U52 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U53 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U54 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U55 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U56 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U57 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U58 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U59 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U60 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U61 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U62 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U63 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U64 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U65 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U66 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U67 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U68 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U69 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U70 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U71 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U72 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U73 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U74 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U75 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U76 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U77 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U78 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U79 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U80 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U81 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U82 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U83 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U84 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U85 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U86 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U87 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U88 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U89 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U90 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U91 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U92 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U93 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U94 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U95 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U96 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U97 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U98 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U99 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U100 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U101 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U102 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U103 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U104 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U105 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U106 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U107 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U108 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U109 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U110 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U111 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U112 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U113 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U114 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U115 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U116 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U117 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U118 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U119 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U120 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U121 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U122 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U123 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U124 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U125 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U126 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U127 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
endmodule


module BWAdder_39 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U3 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U4 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U5 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U6 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U7 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U8 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U9 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U10 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U11 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U12 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U13 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U14 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U15 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U16 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U17 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U18 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U19 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U20 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U21 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U22 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U23 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U24 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U25 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U26 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U27 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U28 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U29 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U30 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U31 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U32 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U33 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U34 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U35 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U36 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U37 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U38 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U39 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U40 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U41 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U42 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U43 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U44 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U45 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U46 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U47 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U48 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U49 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U50 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U51 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U52 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U53 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U54 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U55 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U56 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U57 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U58 ( .A(n59), .ZN(carry[63]) );
  INV_X1 U59 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U60 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U61 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U62 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U63 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U64 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U65 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U66 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U67 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U68 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U69 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U70 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U71 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U72 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U73 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U74 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  AOI22_X1 U75 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U76 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U77 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U78 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U79 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U80 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U81 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U82 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U83 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U84 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U85 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U86 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U87 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U88 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U89 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U90 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U91 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U92 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U93 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U94 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U95 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U96 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U97 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U98 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U99 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U100 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U101 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U102 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U103 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U104 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U105 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U106 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U107 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U108 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U109 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U110 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U111 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U112 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U113 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U114 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U115 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U116 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U117 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U118 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U119 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U120 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U121 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U122 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U123 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U124 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U125 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U126 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U127 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
endmodule


module BWAdder_40 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199;
  assign carry[0] = 1'b0;

  XOR2_X1 U129 ( .A(c[8]), .B(n198), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n197), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n196), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n195), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n195) );
  XOR2_X1 U134 ( .A(c[62]), .B(n194), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n193), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n192), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n191), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n190), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n189), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n188), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n187), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n186), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n185), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n184), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n183), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n182), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n181), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n180), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n179), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n178), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n177), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n176), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n175), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n174), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n173), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n172), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n171), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n170), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n169), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n168), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n167), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n166), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n165), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n164), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n163), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n162), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n161), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n160), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n159), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n158), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n157), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n156), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n155), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n154), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n153), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n152), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n151), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n150), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n149), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n148), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n147), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n146), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n145), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n144), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n143), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n142), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n141), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n140), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n139), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n138), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n137), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n136), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n198) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n197) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n196) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n191) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n194) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n193) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n192) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n190) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n180) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n189) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n188) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n187) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n186) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n185) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n184) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n183) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n182) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n181) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n179) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n169) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n178) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n177) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n176) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n175) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n174) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n173) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n172) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n171) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n170) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n168) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n158) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n167) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n166) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n165) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n164) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n163) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n162) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n161) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n160) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n159) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n157) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n147) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n156) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n155) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n154) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n153) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n152) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n151) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n150) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n149) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n148) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n146) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n136) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n145) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n144) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n143) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n142) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n141) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n140) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n139) );
  INV_X1 U2 ( .A(c[9]), .ZN(n3) );
  INV_X1 U3 ( .A(b[10]), .ZN(n1) );
  INV_X1 U4 ( .A(b[11]), .ZN(n2) );
  INV_X1 U5 ( .A(b[9]), .ZN(n4) );
  XNOR2_X1 U6 ( .A(a[10]), .B(n1), .ZN(n137) );
  XNOR2_X1 U7 ( .A(a[11]), .B(n2), .ZN(n138) );
  XNOR2_X1 U8 ( .A(n3), .B(n199), .ZN(result[9]) );
  XNOR2_X1 U9 ( .A(a[9]), .B(n4), .ZN(n199) );
  INV_X1 U10 ( .A(n14), .ZN(carry[19]) );
  AOI22_X1 U11 ( .A1(b[18]), .A2(a[18]), .B1(n145), .B2(c[18]), .ZN(n14) );
  INV_X1 U12 ( .A(n16), .ZN(carry[20]) );
  AOI22_X1 U13 ( .A1(b[19]), .A2(a[19]), .B1(n146), .B2(c[19]), .ZN(n16) );
  INV_X1 U14 ( .A(n13), .ZN(carry[18]) );
  AOI22_X1 U15 ( .A1(b[17]), .A2(a[17]), .B1(n144), .B2(c[17]), .ZN(n13) );
  INV_X1 U16 ( .A(n17), .ZN(carry[21]) );
  AOI22_X1 U17 ( .A1(b[20]), .A2(a[20]), .B1(n148), .B2(c[20]), .ZN(n17) );
  INV_X1 U18 ( .A(n18), .ZN(carry[22]) );
  AOI22_X1 U19 ( .A1(b[21]), .A2(a[21]), .B1(n149), .B2(c[21]), .ZN(n18) );
  INV_X1 U20 ( .A(n19), .ZN(carry[23]) );
  AOI22_X1 U21 ( .A1(b[22]), .A2(a[22]), .B1(n150), .B2(c[22]), .ZN(n19) );
  INV_X1 U22 ( .A(n20), .ZN(carry[24]) );
  AOI22_X1 U23 ( .A1(b[23]), .A2(a[23]), .B1(n151), .B2(c[23]), .ZN(n20) );
  INV_X1 U24 ( .A(n21), .ZN(carry[25]) );
  AOI22_X1 U25 ( .A1(b[24]), .A2(a[24]), .B1(n152), .B2(c[24]), .ZN(n21) );
  INV_X1 U26 ( .A(n22), .ZN(carry[26]) );
  AOI22_X1 U27 ( .A1(b[25]), .A2(a[25]), .B1(n153), .B2(c[25]), .ZN(n22) );
  INV_X1 U28 ( .A(n23), .ZN(carry[27]) );
  AOI22_X1 U29 ( .A1(b[26]), .A2(a[26]), .B1(n154), .B2(c[26]), .ZN(n23) );
  INV_X1 U30 ( .A(n24), .ZN(carry[28]) );
  AOI22_X1 U31 ( .A1(b[27]), .A2(a[27]), .B1(n155), .B2(c[27]), .ZN(n24) );
  INV_X1 U32 ( .A(n25), .ZN(carry[29]) );
  AOI22_X1 U33 ( .A1(b[28]), .A2(a[28]), .B1(n156), .B2(c[28]), .ZN(n25) );
  INV_X1 U34 ( .A(n33), .ZN(carry[36]) );
  AOI22_X1 U35 ( .A1(b[35]), .A2(a[35]), .B1(n164), .B2(c[35]), .ZN(n33) );
  INV_X1 U36 ( .A(n34), .ZN(carry[37]) );
  AOI22_X1 U37 ( .A1(b[36]), .A2(a[36]), .B1(n165), .B2(c[36]), .ZN(n34) );
  INV_X1 U38 ( .A(n35), .ZN(carry[38]) );
  AOI22_X1 U39 ( .A1(b[37]), .A2(a[37]), .B1(n166), .B2(c[37]), .ZN(n35) );
  INV_X1 U40 ( .A(n36), .ZN(carry[39]) );
  AOI22_X1 U41 ( .A1(b[38]), .A2(a[38]), .B1(n167), .B2(c[38]), .ZN(n36) );
  INV_X1 U42 ( .A(n38), .ZN(carry[40]) );
  AOI22_X1 U43 ( .A1(b[39]), .A2(a[39]), .B1(n168), .B2(c[39]), .ZN(n38) );
  INV_X1 U44 ( .A(n39), .ZN(carry[41]) );
  AOI22_X1 U45 ( .A1(b[40]), .A2(a[40]), .B1(n170), .B2(c[40]), .ZN(n39) );
  INV_X1 U46 ( .A(n40), .ZN(carry[42]) );
  AOI22_X1 U47 ( .A1(b[41]), .A2(a[41]), .B1(n171), .B2(c[41]), .ZN(n40) );
  INV_X1 U48 ( .A(n27), .ZN(carry[30]) );
  AOI22_X1 U49 ( .A1(b[29]), .A2(a[29]), .B1(n157), .B2(c[29]), .ZN(n27) );
  INV_X1 U50 ( .A(n28), .ZN(carry[31]) );
  AOI22_X1 U51 ( .A1(b[30]), .A2(a[30]), .B1(n159), .B2(c[30]), .ZN(n28) );
  INV_X1 U52 ( .A(n29), .ZN(carry[32]) );
  AOI22_X1 U53 ( .A1(b[31]), .A2(a[31]), .B1(n160), .B2(c[31]), .ZN(n29) );
  INV_X1 U54 ( .A(n30), .ZN(carry[33]) );
  AOI22_X1 U55 ( .A1(b[32]), .A2(a[32]), .B1(n161), .B2(c[32]), .ZN(n30) );
  INV_X1 U56 ( .A(n31), .ZN(carry[34]) );
  AOI22_X1 U57 ( .A1(b[33]), .A2(a[33]), .B1(n162), .B2(c[33]), .ZN(n31) );
  INV_X1 U58 ( .A(n32), .ZN(carry[35]) );
  AOI22_X1 U59 ( .A1(b[34]), .A2(a[34]), .B1(n163), .B2(c[34]), .ZN(n32) );
  INV_X1 U60 ( .A(n41), .ZN(carry[43]) );
  AOI22_X1 U61 ( .A1(b[42]), .A2(a[42]), .B1(n172), .B2(c[42]), .ZN(n41) );
  INV_X1 U62 ( .A(n42), .ZN(carry[44]) );
  AOI22_X1 U63 ( .A1(b[43]), .A2(a[43]), .B1(n173), .B2(c[43]), .ZN(n42) );
  INV_X1 U64 ( .A(n43), .ZN(carry[45]) );
  AOI22_X1 U65 ( .A1(b[44]), .A2(a[44]), .B1(n174), .B2(c[44]), .ZN(n43) );
  INV_X1 U66 ( .A(n53), .ZN(carry[54]) );
  AOI22_X1 U67 ( .A1(b[53]), .A2(a[53]), .B1(n184), .B2(c[53]), .ZN(n53) );
  INV_X1 U68 ( .A(n54), .ZN(carry[55]) );
  AOI22_X1 U69 ( .A1(b[54]), .A2(a[54]), .B1(n185), .B2(c[54]), .ZN(n54) );
  INV_X1 U70 ( .A(n55), .ZN(carry[56]) );
  AOI22_X1 U71 ( .A1(b[55]), .A2(a[55]), .B1(n186), .B2(c[55]), .ZN(n55) );
  INV_X1 U72 ( .A(n44), .ZN(carry[46]) );
  AOI22_X1 U73 ( .A1(b[45]), .A2(a[45]), .B1(n175), .B2(c[45]), .ZN(n44) );
  INV_X1 U74 ( .A(n45), .ZN(carry[47]) );
  AOI22_X1 U75 ( .A1(b[46]), .A2(a[46]), .B1(n176), .B2(c[46]), .ZN(n45) );
  INV_X1 U76 ( .A(n46), .ZN(carry[48]) );
  AOI22_X1 U77 ( .A1(b[47]), .A2(a[47]), .B1(n177), .B2(c[47]), .ZN(n46) );
  INV_X1 U78 ( .A(n47), .ZN(carry[49]) );
  AOI22_X1 U79 ( .A1(b[48]), .A2(a[48]), .B1(n178), .B2(c[48]), .ZN(n47) );
  INV_X1 U80 ( .A(n49), .ZN(carry[50]) );
  AOI22_X1 U81 ( .A1(b[49]), .A2(a[49]), .B1(n179), .B2(c[49]), .ZN(n49) );
  INV_X1 U82 ( .A(n50), .ZN(carry[51]) );
  AOI22_X1 U83 ( .A1(b[50]), .A2(a[50]), .B1(n181), .B2(c[50]), .ZN(n50) );
  INV_X1 U84 ( .A(n51), .ZN(carry[52]) );
  AOI22_X1 U85 ( .A1(b[51]), .A2(a[51]), .B1(n182), .B2(c[51]), .ZN(n51) );
  INV_X1 U86 ( .A(n52), .ZN(carry[53]) );
  AOI22_X1 U87 ( .A1(b[52]), .A2(a[52]), .B1(n183), .B2(c[52]), .ZN(n52) );
  INV_X1 U88 ( .A(n56), .ZN(carry[57]) );
  AOI22_X1 U89 ( .A1(b[56]), .A2(a[56]), .B1(n187), .B2(c[56]), .ZN(n56) );
  INV_X1 U90 ( .A(n57), .ZN(carry[58]) );
  AOI22_X1 U91 ( .A1(b[57]), .A2(a[57]), .B1(n188), .B2(c[57]), .ZN(n57) );
  INV_X1 U92 ( .A(n58), .ZN(carry[59]) );
  AOI22_X1 U93 ( .A1(b[58]), .A2(a[58]), .B1(n189), .B2(c[58]), .ZN(n58) );
  INV_X1 U94 ( .A(n60), .ZN(carry[60]) );
  AOI22_X1 U95 ( .A1(b[59]), .A2(a[59]), .B1(n190), .B2(c[59]), .ZN(n60) );
  INV_X1 U96 ( .A(n61), .ZN(carry[61]) );
  AOI22_X1 U97 ( .A1(b[60]), .A2(a[60]), .B1(n192), .B2(c[60]), .ZN(n61) );
  INV_X1 U98 ( .A(n62), .ZN(carry[62]) );
  AOI22_X1 U99 ( .A1(b[61]), .A2(a[61]), .B1(n193), .B2(c[61]), .ZN(n62) );
  INV_X1 U100 ( .A(n63), .ZN(carry[63]) );
  AOI22_X1 U101 ( .A1(b[62]), .A2(a[62]), .B1(n194), .B2(c[62]), .ZN(n63) );
  INV_X1 U102 ( .A(n12), .ZN(carry[17]) );
  AOI22_X1 U103 ( .A1(b[16]), .A2(a[16]), .B1(n143), .B2(c[16]), .ZN(n12) );
  INV_X1 U104 ( .A(n11), .ZN(carry[16]) );
  AOI22_X1 U105 ( .A1(b[15]), .A2(a[15]), .B1(n142), .B2(c[15]), .ZN(n11) );
  INV_X1 U106 ( .A(n10), .ZN(carry[15]) );
  AOI22_X1 U107 ( .A1(b[14]), .A2(a[14]), .B1(n141), .B2(c[14]), .ZN(n10) );
  INV_X1 U108 ( .A(n8), .ZN(carry[13]) );
  AOI22_X1 U109 ( .A1(b[12]), .A2(a[12]), .B1(n139), .B2(c[12]), .ZN(n8) );
  INV_X1 U110 ( .A(n9), .ZN(carry[14]) );
  AOI22_X1 U111 ( .A1(b[13]), .A2(a[13]), .B1(n140), .B2(c[13]), .ZN(n9) );
  INV_X1 U112 ( .A(n5), .ZN(carry[10]) );
  INV_X1 U113 ( .A(n6), .ZN(carry[11]) );
  AOI22_X1 U114 ( .A1(b[10]), .A2(a[10]), .B1(n137), .B2(c[10]), .ZN(n6) );
  INV_X1 U115 ( .A(n7), .ZN(carry[12]) );
  AOI22_X1 U116 ( .A1(b[11]), .A2(a[11]), .B1(n138), .B2(c[11]), .ZN(n7) );
  INV_X1 U117 ( .A(n15), .ZN(carry[1]) );
  AOI22_X1 U118 ( .A1(b[0]), .A2(a[0]), .B1(n136), .B2(c[0]), .ZN(n15) );
  INV_X1 U119 ( .A(n26), .ZN(carry[2]) );
  AOI22_X1 U120 ( .A1(b[1]), .A2(a[1]), .B1(n147), .B2(c[1]), .ZN(n26) );
  INV_X1 U121 ( .A(n37), .ZN(carry[3]) );
  AOI22_X1 U122 ( .A1(b[2]), .A2(a[2]), .B1(n158), .B2(c[2]), .ZN(n37) );
  INV_X1 U123 ( .A(n48), .ZN(carry[4]) );
  AOI22_X1 U124 ( .A1(b[3]), .A2(a[3]), .B1(n169), .B2(c[3]), .ZN(n48) );
  INV_X1 U125 ( .A(n59), .ZN(carry[5]) );
  AOI22_X1 U126 ( .A1(b[4]), .A2(a[4]), .B1(n180), .B2(c[4]), .ZN(n59) );
  INV_X1 U127 ( .A(n132), .ZN(carry[6]) );
  AOI22_X1 U128 ( .A1(b[5]), .A2(a[5]), .B1(n191), .B2(c[5]), .ZN(n132) );
  INV_X1 U253 ( .A(n135), .ZN(carry[9]) );
  AOI22_X1 U254 ( .A1(b[8]), .A2(a[8]), .B1(n198), .B2(c[8]), .ZN(n135) );
  INV_X1 U255 ( .A(n133), .ZN(carry[7]) );
  AOI22_X1 U256 ( .A1(b[6]), .A2(a[6]), .B1(n196), .B2(c[6]), .ZN(n133) );
  INV_X1 U257 ( .A(n134), .ZN(carry[8]) );
  AOI22_X1 U258 ( .A1(b[7]), .A2(a[7]), .B1(n197), .B2(c[7]), .ZN(n134) );
  AOI22_X1 U259 ( .A1(b[9]), .A2(a[9]), .B1(n199), .B2(c[9]), .ZN(n5) );
endmodule


module BWAdder_41 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n65, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(n204), .B(c[9]), .Z(result[9]) );
  XOR2_X1 U129 ( .A(n7), .B(c[8]), .Z(result[8]) );
  XOR2_X1 U130 ( .A(n203), .B(c[7]), .Z(result[7]) );
  XOR2_X1 U131 ( .A(n202), .B(c[6]), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n201), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n201) );
  XOR2_X1 U134 ( .A(c[62]), .B(n200), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n199), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n198), .Z(result[60]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n196), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n195), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n194), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n193), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n192), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n191), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n190), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n189), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n188), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n187), .Z(result[50]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n185), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n184), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n183), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n182), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n181), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n180), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n179), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n178), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n177), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n176), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n175), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n174), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n173), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n172), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n171), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n170), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n169), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n168), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n167), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n166), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n165), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n164), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n163), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n162), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n161), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n160), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n159), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n158), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n157), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n156), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n155), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n154), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n153), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n152), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n151), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n150), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n149), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n148), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n147), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n146), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n145), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n144), .Z(result[11]) );
  XOR2_X1 U191 ( .A(n143), .B(c[10]), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n142), .Z(result[0]) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n203) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n202) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n197) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n200) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n199) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n198) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n196) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n186) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n195) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n194) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n193) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n192) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n191) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n190) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n189) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n188) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n187) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n185) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n175) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n184) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n183) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n182) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n181) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n180) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n179) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n178) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n177) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n176) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n174) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n164) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n173) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n172) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n171) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n170) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n169) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n168) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n167) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n166) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n165) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n163) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n153) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n162) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n161) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n160) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n159) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n158) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n157) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n156) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n155) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n154) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n152) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n142) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n151) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n150) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n149) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n148) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n147) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n146) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n145) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n144) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n143) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n204) );
  CLKBUF_X1 U2 ( .A(a[6]), .Z(n1) );
  INV_X1 U3 ( .A(c[4]), .ZN(n5) );
  INV_X1 U4 ( .A(c[5]), .ZN(n6) );
  CLKBUF_X1 U5 ( .A(b[7]), .Z(n2) );
  CLKBUF_X1 U6 ( .A(a[8]), .Z(n3) );
  CLKBUF_X1 U7 ( .A(b[4]), .Z(n4) );
  XNOR2_X1 U8 ( .A(n5), .B(n186), .ZN(result[4]) );
  XNOR2_X1 U9 ( .A(n197), .B(n6), .ZN(result[5]) );
  XOR2_X1 U10 ( .A(a[8]), .B(b[8]), .Z(n7) );
  INV_X1 U11 ( .A(n141), .ZN(carry[9]) );
  INV_X1 U12 ( .A(n9), .ZN(carry[10]) );
  INV_X1 U13 ( .A(n10), .ZN(carry[11]) );
  INV_X1 U14 ( .A(n11), .ZN(carry[12]) );
  AOI22_X1 U15 ( .A1(b[11]), .A2(a[11]), .B1(n144), .B2(c[11]), .ZN(n11) );
  INV_X1 U16 ( .A(n22), .ZN(carry[22]) );
  AOI22_X1 U17 ( .A1(b[21]), .A2(a[21]), .B1(n155), .B2(c[21]), .ZN(n22) );
  INV_X1 U18 ( .A(n21), .ZN(carry[21]) );
  AOI22_X1 U19 ( .A1(b[20]), .A2(a[20]), .B1(n154), .B2(c[20]), .ZN(n21) );
  INV_X1 U20 ( .A(n12), .ZN(carry[13]) );
  AOI22_X1 U21 ( .A1(b[12]), .A2(a[12]), .B1(n145), .B2(c[12]), .ZN(n12) );
  INV_X1 U22 ( .A(n20), .ZN(carry[20]) );
  AOI22_X1 U23 ( .A1(b[19]), .A2(a[19]), .B1(n152), .B2(c[19]), .ZN(n20) );
  INV_X1 U24 ( .A(n16), .ZN(carry[17]) );
  AOI22_X1 U25 ( .A1(b[16]), .A2(a[16]), .B1(n149), .B2(c[16]), .ZN(n16) );
  INV_X1 U26 ( .A(n13), .ZN(carry[14]) );
  AOI22_X1 U27 ( .A1(b[13]), .A2(a[13]), .B1(n146), .B2(c[13]), .ZN(n13) );
  INV_X1 U28 ( .A(n15), .ZN(carry[16]) );
  AOI22_X1 U29 ( .A1(b[15]), .A2(a[15]), .B1(n148), .B2(c[15]), .ZN(n15) );
  INV_X1 U30 ( .A(n14), .ZN(carry[15]) );
  AOI22_X1 U31 ( .A1(b[14]), .A2(a[14]), .B1(n147), .B2(c[14]), .ZN(n14) );
  INV_X1 U32 ( .A(n17), .ZN(carry[18]) );
  AOI22_X1 U33 ( .A1(b[17]), .A2(a[17]), .B1(n150), .B2(c[17]), .ZN(n17) );
  INV_X1 U34 ( .A(n18), .ZN(carry[19]) );
  AOI22_X1 U35 ( .A1(b[18]), .A2(a[18]), .B1(n151), .B2(c[18]), .ZN(n18) );
  INV_X1 U36 ( .A(n23), .ZN(carry[23]) );
  AOI22_X1 U37 ( .A1(b[22]), .A2(a[22]), .B1(n156), .B2(c[22]), .ZN(n23) );
  INV_X1 U38 ( .A(n24), .ZN(carry[24]) );
  AOI22_X1 U39 ( .A1(b[23]), .A2(a[23]), .B1(n157), .B2(c[23]), .ZN(n24) );
  INV_X1 U40 ( .A(n25), .ZN(carry[25]) );
  AOI22_X1 U41 ( .A1(b[24]), .A2(a[24]), .B1(n158), .B2(c[24]), .ZN(n25) );
  INV_X1 U42 ( .A(n26), .ZN(carry[26]) );
  AOI22_X1 U43 ( .A1(b[25]), .A2(a[25]), .B1(n159), .B2(c[25]), .ZN(n26) );
  INV_X1 U44 ( .A(n27), .ZN(carry[27]) );
  AOI22_X1 U45 ( .A1(b[26]), .A2(a[26]), .B1(n160), .B2(c[26]), .ZN(n27) );
  INV_X1 U46 ( .A(n28), .ZN(carry[28]) );
  AOI22_X1 U47 ( .A1(b[27]), .A2(a[27]), .B1(n161), .B2(c[27]), .ZN(n28) );
  INV_X1 U48 ( .A(n29), .ZN(carry[29]) );
  AOI22_X1 U49 ( .A1(b[28]), .A2(a[28]), .B1(n162), .B2(c[28]), .ZN(n29) );
  INV_X1 U50 ( .A(n31), .ZN(carry[30]) );
  AOI22_X1 U51 ( .A1(b[29]), .A2(a[29]), .B1(n163), .B2(c[29]), .ZN(n31) );
  INV_X1 U52 ( .A(n32), .ZN(carry[31]) );
  AOI22_X1 U53 ( .A1(b[30]), .A2(a[30]), .B1(n165), .B2(c[30]), .ZN(n32) );
  INV_X1 U54 ( .A(n33), .ZN(carry[32]) );
  AOI22_X1 U55 ( .A1(b[31]), .A2(a[31]), .B1(n166), .B2(c[31]), .ZN(n33) );
  INV_X1 U56 ( .A(n34), .ZN(carry[33]) );
  AOI22_X1 U57 ( .A1(b[32]), .A2(a[32]), .B1(n167), .B2(c[32]), .ZN(n34) );
  INV_X1 U58 ( .A(n37), .ZN(carry[36]) );
  AOI22_X1 U59 ( .A1(b[35]), .A2(a[35]), .B1(n170), .B2(c[35]), .ZN(n37) );
  INV_X1 U60 ( .A(n38), .ZN(carry[37]) );
  AOI22_X1 U61 ( .A1(b[36]), .A2(a[36]), .B1(n171), .B2(c[36]), .ZN(n38) );
  INV_X1 U62 ( .A(n39), .ZN(carry[38]) );
  AOI22_X1 U63 ( .A1(b[37]), .A2(a[37]), .B1(n172), .B2(c[37]), .ZN(n39) );
  INV_X1 U64 ( .A(n40), .ZN(carry[39]) );
  AOI22_X1 U65 ( .A1(b[38]), .A2(a[38]), .B1(n173), .B2(c[38]), .ZN(n40) );
  INV_X1 U66 ( .A(n42), .ZN(carry[40]) );
  AOI22_X1 U67 ( .A1(b[39]), .A2(a[39]), .B1(n174), .B2(c[39]), .ZN(n42) );
  INV_X1 U68 ( .A(n43), .ZN(carry[41]) );
  AOI22_X1 U69 ( .A1(b[40]), .A2(a[40]), .B1(n176), .B2(c[40]), .ZN(n43) );
  INV_X1 U70 ( .A(n44), .ZN(carry[42]) );
  AOI22_X1 U71 ( .A1(b[41]), .A2(a[41]), .B1(n177), .B2(c[41]), .ZN(n44) );
  INV_X1 U72 ( .A(n45), .ZN(carry[43]) );
  AOI22_X1 U73 ( .A1(b[42]), .A2(a[42]), .B1(n178), .B2(c[42]), .ZN(n45) );
  INV_X1 U74 ( .A(n35), .ZN(carry[34]) );
  AOI22_X1 U75 ( .A1(b[33]), .A2(a[33]), .B1(n168), .B2(c[33]), .ZN(n35) );
  INV_X1 U76 ( .A(n36), .ZN(carry[35]) );
  AOI22_X1 U77 ( .A1(b[34]), .A2(a[34]), .B1(n169), .B2(c[34]), .ZN(n36) );
  INV_X1 U78 ( .A(n59), .ZN(carry[56]) );
  AOI22_X1 U79 ( .A1(b[55]), .A2(a[55]), .B1(n192), .B2(c[55]), .ZN(n59) );
  INV_X1 U80 ( .A(n46), .ZN(carry[44]) );
  AOI22_X1 U81 ( .A1(b[43]), .A2(a[43]), .B1(n179), .B2(c[43]), .ZN(n46) );
  INV_X1 U82 ( .A(n47), .ZN(carry[45]) );
  AOI22_X1 U83 ( .A1(b[44]), .A2(a[44]), .B1(n180), .B2(c[44]), .ZN(n47) );
  INV_X1 U84 ( .A(n48), .ZN(carry[46]) );
  AOI22_X1 U85 ( .A1(b[45]), .A2(a[45]), .B1(n181), .B2(c[45]), .ZN(n48) );
  INV_X1 U86 ( .A(n49), .ZN(carry[47]) );
  AOI22_X1 U87 ( .A1(b[46]), .A2(a[46]), .B1(n182), .B2(c[46]), .ZN(n49) );
  INV_X1 U88 ( .A(n50), .ZN(carry[48]) );
  AOI22_X1 U89 ( .A1(b[47]), .A2(a[47]), .B1(n183), .B2(c[47]), .ZN(n50) );
  INV_X1 U90 ( .A(n51), .ZN(carry[49]) );
  AOI22_X1 U91 ( .A1(b[48]), .A2(a[48]), .B1(n184), .B2(c[48]), .ZN(n51) );
  INV_X1 U92 ( .A(n53), .ZN(carry[50]) );
  AOI22_X1 U93 ( .A1(b[49]), .A2(a[49]), .B1(n185), .B2(c[49]), .ZN(n53) );
  INV_X1 U94 ( .A(n54), .ZN(carry[51]) );
  AOI22_X1 U95 ( .A1(b[50]), .A2(a[50]), .B1(n187), .B2(c[50]), .ZN(n54) );
  INV_X1 U96 ( .A(n55), .ZN(carry[52]) );
  AOI22_X1 U97 ( .A1(b[51]), .A2(a[51]), .B1(n188), .B2(c[51]), .ZN(n55) );
  INV_X1 U98 ( .A(n56), .ZN(carry[53]) );
  AOI22_X1 U99 ( .A1(b[52]), .A2(a[52]), .B1(n189), .B2(c[52]), .ZN(n56) );
  INV_X1 U100 ( .A(n57), .ZN(carry[54]) );
  AOI22_X1 U101 ( .A1(b[53]), .A2(a[53]), .B1(n190), .B2(c[53]), .ZN(n57) );
  INV_X1 U102 ( .A(n58), .ZN(carry[55]) );
  AOI22_X1 U103 ( .A1(b[54]), .A2(a[54]), .B1(n191), .B2(c[54]), .ZN(n58) );
  INV_X1 U104 ( .A(n60), .ZN(carry[57]) );
  AOI22_X1 U105 ( .A1(b[56]), .A2(a[56]), .B1(n193), .B2(c[56]), .ZN(n60) );
  INV_X1 U106 ( .A(n61), .ZN(carry[58]) );
  AOI22_X1 U107 ( .A1(b[57]), .A2(a[57]), .B1(n194), .B2(c[57]), .ZN(n61) );
  INV_X1 U108 ( .A(n62), .ZN(carry[59]) );
  AOI22_X1 U109 ( .A1(b[58]), .A2(a[58]), .B1(n195), .B2(c[58]), .ZN(n62) );
  INV_X1 U110 ( .A(n65), .ZN(carry[60]) );
  AOI22_X1 U111 ( .A1(b[59]), .A2(a[59]), .B1(n196), .B2(c[59]), .ZN(n65) );
  INV_X1 U112 ( .A(n135), .ZN(carry[61]) );
  AOI22_X1 U113 ( .A1(b[60]), .A2(a[60]), .B1(n198), .B2(c[60]), .ZN(n135) );
  INV_X1 U114 ( .A(n136), .ZN(carry[62]) );
  AOI22_X1 U115 ( .A1(b[61]), .A2(a[61]), .B1(n199), .B2(c[61]), .ZN(n136) );
  INV_X1 U116 ( .A(n137), .ZN(carry[63]) );
  AOI22_X1 U117 ( .A1(b[62]), .A2(a[62]), .B1(n200), .B2(c[62]), .ZN(n137) );
  INV_X1 U118 ( .A(n138), .ZN(carry[6]) );
  INV_X1 U119 ( .A(n63), .ZN(carry[5]) );
  INV_X1 U120 ( .A(n52), .ZN(carry[4]) );
  INV_X1 U121 ( .A(n140), .ZN(carry[8]) );
  INV_X1 U122 ( .A(n19), .ZN(carry[1]) );
  AOI22_X1 U123 ( .A1(b[0]), .A2(a[0]), .B1(n142), .B2(c[0]), .ZN(n19) );
  INV_X1 U124 ( .A(n30), .ZN(carry[2]) );
  AOI22_X1 U125 ( .A1(b[1]), .A2(a[1]), .B1(n153), .B2(c[1]), .ZN(n30) );
  INV_X1 U126 ( .A(n41), .ZN(carry[3]) );
  AOI22_X1 U127 ( .A1(b[2]), .A2(a[2]), .B1(n164), .B2(c[2]), .ZN(n41) );
  CLKBUF_X1 U137 ( .A(b[6]), .Z(n8) );
  AOI22_X1 U148 ( .A1(b[3]), .A2(a[3]), .B1(n175), .B2(c[3]), .ZN(n52) );
  AOI22_X1 U193 ( .A1(b[10]), .A2(a[10]), .B1(n143), .B2(c[10]), .ZN(n10) );
  INV_X1 U256 ( .A(n139), .ZN(carry[7]) );
  AOI22_X1 U257 ( .A1(b[9]), .A2(a[9]), .B1(n204), .B2(c[9]), .ZN(n9) );
  AOI22_X1 U258 ( .A1(n4), .A2(a[4]), .B1(n186), .B2(c[4]), .ZN(n63) );
  AOI22_X1 U259 ( .A1(n8), .A2(n1), .B1(n202), .B2(c[6]), .ZN(n139) );
  AOI22_X1 U260 ( .A1(b[5]), .A2(a[5]), .B1(n197), .B2(c[5]), .ZN(n138) );
  AOI22_X1 U261 ( .A1(n2), .A2(a[7]), .B1(n203), .B2(c[7]), .ZN(n140) );
  AOI22_X1 U262 ( .A1(b[8]), .A2(n3), .B1(n7), .B2(c[8]), .ZN(n141) );
endmodule


module BWAdder_42 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U3 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U4 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U5 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U6 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U7 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U8 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U9 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U10 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U11 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U12 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U13 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U14 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U15 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U16 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U17 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U18 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U19 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U20 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U21 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U22 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U23 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U24 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U25 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U26 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U27 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U28 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U29 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U30 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U31 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U32 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U33 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U34 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U35 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U36 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U37 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U38 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U39 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U40 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U41 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U42 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U43 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U44 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U45 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U46 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U47 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U48 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U49 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U50 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U51 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U52 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U53 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U54 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U55 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U56 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U57 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U58 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U59 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U60 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U61 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U62 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U63 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U64 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U65 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U66 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U67 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U68 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U69 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U70 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U71 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U72 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U73 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U74 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U75 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U76 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U77 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U78 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U79 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U80 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U81 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U82 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U83 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U84 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U85 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U86 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U87 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U88 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U89 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U90 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U91 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U92 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U93 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U94 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U95 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U96 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U97 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U98 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U99 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U100 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U101 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U102 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U103 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U104 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U105 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U106 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U107 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U108 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U109 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U110 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U111 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U112 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U113 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U114 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U115 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U116 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U117 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U118 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U119 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U120 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U121 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U122 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U123 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U124 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U125 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U126 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U127 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
endmodule


module BWAdder_43 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U3 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U4 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U5 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U6 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U7 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U8 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U9 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U10 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U11 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U12 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U13 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U14 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U15 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U16 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U17 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U18 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U19 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U20 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U21 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U22 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U23 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U24 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U25 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U26 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U27 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U28 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U29 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U30 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U31 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U32 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U33 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U34 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U35 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U36 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U37 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U38 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U39 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U40 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U41 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U42 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U43 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U44 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U45 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U46 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U47 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U48 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U49 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U50 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U51 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U52 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U53 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U54 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U55 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U56 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U57 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U58 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U59 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U60 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U61 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U62 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U63 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U64 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U65 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U66 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U67 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U68 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U69 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U70 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U71 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U72 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U73 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U74 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U75 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U76 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U77 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U78 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U79 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U80 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U81 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U82 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U83 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U84 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U85 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U86 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U87 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U88 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U89 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U90 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U91 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U92 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U93 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U94 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U95 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U96 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U97 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U98 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U99 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U100 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U101 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U102 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U103 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U104 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U105 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U106 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U107 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U108 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U109 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U110 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U111 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U112 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U113 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U114 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U115 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U116 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U117 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U118 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U119 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U120 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U121 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U122 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U123 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U124 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U125 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U126 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U127 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
endmodule


module BWAdder_44 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U3 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U4 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U5 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U6 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U7 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U8 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U9 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U10 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U11 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U12 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U13 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U14 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U15 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U16 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U17 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U18 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U19 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U20 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U21 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U22 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U23 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U24 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U25 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U26 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U27 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U28 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U29 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U30 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U31 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U32 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U33 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U34 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U35 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U36 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U37 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U38 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U39 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U40 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U41 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U42 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U43 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U44 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U45 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U46 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U47 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U48 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U49 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U50 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U51 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U52 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U53 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U54 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U55 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U56 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U57 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U58 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U59 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U60 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U61 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U62 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U63 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U64 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U65 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U66 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U67 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U68 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U69 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U70 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U71 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U72 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U73 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U74 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U75 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U76 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U77 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U78 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U79 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U80 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U81 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U82 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U83 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U84 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U85 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U86 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U87 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U88 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U89 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U90 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U91 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U92 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U93 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U94 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U95 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U96 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U97 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U98 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U99 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U100 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U101 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U102 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U103 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U104 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U105 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U106 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U107 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U108 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U109 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U110 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U111 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U112 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U113 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U114 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U115 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U116 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U117 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U118 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U120 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U121 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U122 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U123 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U124 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U125 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U126 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U127 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
endmodule


module BWAdder_45 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U3 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U4 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U5 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U6 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U7 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U8 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U9 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U10 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U11 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U12 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U13 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U14 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U15 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U16 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U17 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U18 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U19 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U20 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U21 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U22 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U23 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U24 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U25 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U26 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U27 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U28 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U29 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U30 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U31 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U32 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U33 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U34 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U35 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U36 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U37 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U38 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U39 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U40 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U41 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U42 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U43 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U44 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U45 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U46 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U47 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U48 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U49 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U50 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U51 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U52 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U53 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U54 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U55 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U56 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U57 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U58 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U59 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U60 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U61 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U62 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U63 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U64 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U65 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U66 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U67 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U68 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U69 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U70 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U71 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U72 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U73 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U74 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U75 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U76 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U77 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U78 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U79 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U80 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U81 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U82 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U83 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U84 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U85 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U86 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U87 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U88 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U89 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U90 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U91 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U92 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U93 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U94 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U95 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U96 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U97 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U98 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U99 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U100 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U101 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U102 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U103 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U104 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U105 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U106 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U107 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U108 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U109 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U110 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U111 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U112 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U113 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U114 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U115 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U116 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U117 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U118 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U119 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U120 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U121 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U122 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U123 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U124 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U125 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U126 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U127 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
endmodule


module BWAdder_46 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U3 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U4 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U5 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U6 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U7 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U8 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U9 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U10 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U11 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U12 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U13 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U14 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U15 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U16 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U17 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U18 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U19 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U20 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U21 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U22 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U23 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U24 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U25 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U26 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U27 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U28 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U29 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U30 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U31 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U32 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U33 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U34 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U35 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U36 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U37 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U38 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U39 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U40 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U41 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U42 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U43 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U44 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U45 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U46 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U47 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U48 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U49 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U50 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U51 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U52 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U53 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U54 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U55 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U56 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U57 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U58 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U59 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U60 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U61 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U62 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U63 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U64 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U65 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U66 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U67 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U68 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U69 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U70 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U71 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U72 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U73 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U74 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U75 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U76 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U77 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U78 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U79 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U80 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U81 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U82 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U83 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U84 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U85 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U86 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U87 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U88 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U89 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U90 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U91 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U92 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U93 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U94 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U95 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U96 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U97 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U98 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U99 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U100 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U101 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U102 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U103 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U104 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U105 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U106 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U107 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U108 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U109 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U110 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U111 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U112 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U113 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U114 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U115 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U116 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U117 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U118 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U119 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U120 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U121 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U122 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U123 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U124 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U125 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U126 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U127 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
endmodule


module BWAdder_47 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U3 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U4 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U5 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U6 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U7 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U8 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U9 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U10 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U11 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U12 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U13 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U14 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U15 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U16 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U17 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U18 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U19 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U20 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U21 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U22 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U23 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U24 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U25 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U26 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U27 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U28 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U29 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U30 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U31 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U32 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U33 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U34 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U35 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U36 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U37 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U38 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U39 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U40 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U41 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U42 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U43 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U44 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U45 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U46 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U47 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U48 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U49 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U50 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U51 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U52 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U53 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U54 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U55 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U56 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U57 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U58 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U59 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U60 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U61 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U62 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U63 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U64 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U65 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U66 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U67 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U68 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U69 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U70 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U71 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U72 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U73 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U74 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U75 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U76 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U77 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U78 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U79 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U80 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U81 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U82 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U83 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U84 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U85 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U86 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U87 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U88 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U89 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U90 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U91 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U92 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U93 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U94 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U95 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U96 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U97 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U98 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U99 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U100 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U101 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U102 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U103 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U104 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U105 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U106 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U107 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U108 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U109 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U110 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U111 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U112 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U113 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U114 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U115 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U116 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U117 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U118 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U119 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U120 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U121 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U122 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U123 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U124 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U125 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U126 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U127 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
endmodule


module BWAdder_48 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U3 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U4 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U5 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U6 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U7 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U8 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U9 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U10 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U11 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U12 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U13 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U14 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U15 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U16 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U17 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U18 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U19 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U20 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U21 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U22 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U23 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U24 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U25 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U26 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U27 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U28 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U29 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U30 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U31 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U32 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U33 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U34 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U35 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U36 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U37 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  AOI22_X1 U38 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U39 ( .A(n59), .ZN(carry[63]) );
  INV_X1 U40 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U41 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U42 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U43 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U44 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U45 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U46 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U47 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U48 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U49 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U50 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U51 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U52 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U53 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U54 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U55 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U56 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U57 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U58 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U59 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U60 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U61 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U62 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U63 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U64 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U65 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U66 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U67 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U68 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U69 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U70 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U71 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U72 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U73 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U74 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U75 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U76 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U77 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U78 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U79 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U80 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U81 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U82 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U83 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U84 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U85 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U86 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U87 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U88 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U89 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U90 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U91 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U92 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U93 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U94 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U95 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U96 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U97 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U98 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U99 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U100 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U101 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U102 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U103 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U104 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U105 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U106 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U107 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U108 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U109 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U110 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U111 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U112 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U113 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U114 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U115 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U116 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U117 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U118 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U119 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U120 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U121 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U122 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U123 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U124 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U125 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U126 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U127 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
endmodule


module BWAdder_49 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U3 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U4 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U5 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U6 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U7 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U8 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U9 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U10 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U11 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U12 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U13 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U14 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U15 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U16 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U17 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U18 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U19 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U20 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U21 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U22 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U23 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U24 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U25 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U26 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U27 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U28 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U29 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U30 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U31 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U32 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U33 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U34 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U35 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U36 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U37 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U38 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U39 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U40 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U41 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U42 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U43 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U44 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U45 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U46 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U47 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U48 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U49 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U50 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U51 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U52 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U53 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U54 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U55 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U56 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U57 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U58 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U59 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U60 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U61 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U62 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U63 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U64 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U65 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U66 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U67 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U68 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U69 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U70 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U71 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U72 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U73 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U74 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U75 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U76 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U77 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U78 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U79 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U80 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U81 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U82 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U83 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U84 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U85 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U86 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U87 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U88 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U89 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U90 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U91 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U92 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U93 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U94 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U95 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U96 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U97 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U98 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U99 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U100 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U101 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U102 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U103 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U104 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U105 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U106 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U107 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U108 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U109 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U110 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U111 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U112 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U113 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U114 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U115 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U116 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U117 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U118 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U119 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U120 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U121 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U122 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U123 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U124 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U125 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U126 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U127 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
endmodule


module BWAdder_50 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U3 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U4 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U5 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U6 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U7 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U8 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U9 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U10 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U11 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U12 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U13 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U14 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U15 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U16 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U17 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U18 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U19 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U20 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U21 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U22 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U23 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U24 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U25 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U26 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U27 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U28 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U29 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U30 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U31 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U32 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U33 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U34 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U35 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U36 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U37 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U38 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U39 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U40 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U41 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U42 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U43 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U44 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U45 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U46 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U47 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U48 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U49 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U50 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U51 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U52 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U53 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U54 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U55 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U56 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U57 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U58 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U59 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U60 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U61 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U62 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U63 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U64 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U65 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U66 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U67 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U68 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U69 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U70 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U71 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U72 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U73 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U74 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U75 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U76 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U77 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U78 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U79 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U80 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U81 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U82 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U83 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U84 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U85 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U86 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U87 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U88 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U89 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U90 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U91 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U92 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U93 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U94 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U95 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U96 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U97 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U98 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U99 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U100 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U101 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U102 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U103 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U104 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U105 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U106 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U107 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U108 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U109 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U110 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U111 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U112 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U113 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U114 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U115 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U116 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U117 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U118 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U119 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U120 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U121 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U122 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U123 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U124 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U125 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U126 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U127 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
endmodule


module BWAdder_51 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U3 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U4 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U5 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U6 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U7 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U8 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U9 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U10 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U11 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U12 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U13 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U14 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U15 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U16 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U17 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U18 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U19 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U20 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U21 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U22 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U23 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U24 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U25 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U26 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U27 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U28 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U29 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U30 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U31 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U32 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U33 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U34 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U35 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U36 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U37 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U38 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U39 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U40 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U41 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U42 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U43 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U44 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U45 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U46 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U47 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U48 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U49 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U50 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U51 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U52 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U53 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U54 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U55 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U56 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U57 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U58 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U59 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U60 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U61 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U62 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U63 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U64 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U65 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U66 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U67 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U68 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U69 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U70 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U71 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U72 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U73 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U74 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U75 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U76 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U77 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U78 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U79 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U80 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U81 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U82 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U83 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U84 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U85 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U86 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U87 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U88 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U89 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U90 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U91 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U92 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U93 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U94 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U95 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U96 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U97 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U98 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U99 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U100 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U101 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U102 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U103 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U104 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U105 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U106 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U107 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U108 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U109 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U110 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U111 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U112 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U113 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U114 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U115 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U116 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U117 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U118 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U119 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U120 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U121 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U122 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U123 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U124 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U125 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U126 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U127 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
endmodule


module BWAdder_52 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U3 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U4 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U5 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U6 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U7 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U8 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U9 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U10 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U11 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U12 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U13 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U14 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U15 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U16 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U17 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U18 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U19 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U20 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U21 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U22 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U23 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U24 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U25 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U26 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U27 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U28 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U29 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U30 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U31 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U32 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U33 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U34 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U35 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U36 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U37 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U38 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U39 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U40 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U41 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U42 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U43 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U44 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U45 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U46 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U47 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U48 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U49 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U50 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U51 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U52 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U53 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U54 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U55 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U56 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U57 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U58 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U59 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U60 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U61 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U62 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U63 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U64 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U65 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U66 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U67 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U68 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U69 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U70 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U71 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U72 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U73 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U74 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U75 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U76 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U78 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U79 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U80 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U81 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U82 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U83 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U84 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U85 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U86 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U87 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U88 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U89 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U90 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U91 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U92 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U93 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U94 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U95 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U96 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U97 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U98 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U99 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U100 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U101 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U102 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U103 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U104 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U105 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U106 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U107 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U108 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U109 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U110 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U111 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U112 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U113 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U114 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U115 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U116 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U117 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U118 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U119 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U120 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U121 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U122 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U123 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U124 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U125 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U126 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U127 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
endmodule


module BWAdder_53 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U3 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U4 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U5 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U6 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U7 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U8 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U9 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U10 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U11 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U12 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U13 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U14 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U15 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U16 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U17 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U18 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U19 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U20 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U21 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U22 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U23 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U24 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U25 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U26 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U27 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U28 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U29 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U30 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U31 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U32 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U33 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U34 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U35 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U36 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U37 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U38 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U39 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U40 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U41 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U42 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U43 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U44 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U45 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U46 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U47 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U48 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U49 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U50 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U51 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U52 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U53 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U54 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U55 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U56 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U57 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U58 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U59 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U60 ( .A(n59), .ZN(carry[63]) );
  INV_X1 U61 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U62 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U63 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U64 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U65 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U66 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U67 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U68 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  AOI22_X1 U69 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U70 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U71 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U72 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U73 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U74 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U75 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U76 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U77 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U78 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U79 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U80 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U81 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U82 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U83 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U84 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U85 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U86 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U87 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U88 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U89 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U90 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U91 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U92 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U93 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U94 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U95 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U96 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U97 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U98 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U99 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U100 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U101 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U102 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U103 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U104 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U105 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U106 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U107 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U108 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U109 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U110 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U111 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U112 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U113 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U114 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U115 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U116 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U117 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U118 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U119 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U120 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U121 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U122 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U123 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U124 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U125 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U126 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U127 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
endmodule


module BWAdder_54 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U3 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U4 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U5 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U6 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U7 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U8 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U9 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U10 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U11 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U12 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U13 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U14 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U15 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U16 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U17 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U18 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U19 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U20 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U21 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U22 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U23 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U24 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U25 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U26 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U27 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U28 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U29 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U30 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U31 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U32 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U33 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U34 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U35 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U36 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U37 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U38 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U39 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U40 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U41 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U42 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U43 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U44 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U45 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U46 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U47 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U48 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U49 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U50 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U51 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U52 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U53 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U54 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U55 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U56 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U57 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U58 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U59 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U60 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U61 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U62 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U63 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U64 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U65 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U66 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U67 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U68 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U69 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U70 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U71 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U72 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U73 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U74 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U75 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U76 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U77 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U78 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U79 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U80 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U81 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U82 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U83 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U84 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U85 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U86 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U87 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U88 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U89 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U90 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U91 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U92 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U93 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U94 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U95 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U96 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U97 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U98 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U99 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U100 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U101 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U102 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U103 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U104 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U105 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U106 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U107 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U108 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U109 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U110 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U111 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U112 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U113 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U114 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U115 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U116 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U117 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U118 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U119 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U120 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U121 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U122 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U123 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U124 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U125 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U126 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U127 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
endmodule


module BWAdder_55 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U3 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U4 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U5 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U6 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U7 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U8 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U9 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U10 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U11 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U12 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U13 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U14 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U15 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U16 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U17 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U18 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U19 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U20 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U21 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U22 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U23 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U24 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U25 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U26 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U27 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U28 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U29 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U30 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U31 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U32 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U33 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U34 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U35 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U36 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U37 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U38 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U39 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U40 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U41 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U42 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U43 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U44 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U45 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U46 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U47 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U48 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U49 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U50 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U51 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U52 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U53 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U54 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U55 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U56 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U57 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U58 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U59 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U60 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U61 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U62 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U63 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U64 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U65 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U66 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U67 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U68 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U69 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U70 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U71 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U72 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U73 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U74 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U75 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U76 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U77 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U78 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U79 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U80 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U81 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U82 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U83 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U84 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U85 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U86 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U87 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U88 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U89 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U90 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U91 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U92 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U93 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U94 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U95 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U96 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U97 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U98 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U99 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U100 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U101 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U102 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U103 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U104 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U105 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U106 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U107 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U108 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U109 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U110 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U111 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U112 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U113 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U114 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U115 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U116 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U117 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U118 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U119 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U120 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U121 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U122 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U123 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U124 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U125 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U126 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U127 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
endmodule


module BWAdder_56 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U3 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U4 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U5 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U6 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U7 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U8 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U9 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U10 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U11 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U12 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U13 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U14 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U15 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U16 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U17 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U18 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U19 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U20 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U21 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U22 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U23 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U24 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U25 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U26 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U27 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U28 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U29 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U30 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U31 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U32 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U33 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U34 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U35 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U36 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U37 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U38 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U39 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U40 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U41 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U42 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U43 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U44 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U45 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U46 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U47 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U48 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U49 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U50 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U51 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U52 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U53 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U54 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U55 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U56 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U57 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U58 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U59 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U60 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U61 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U62 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U63 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U64 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U65 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U66 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U67 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U68 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U69 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U70 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U71 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U72 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U73 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U74 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U75 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U76 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U77 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U78 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U79 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U80 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U81 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U82 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U83 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U84 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U85 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U86 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U87 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U88 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U89 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U90 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U91 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U92 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U93 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U94 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U95 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U96 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U97 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U98 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U99 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U100 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U101 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U102 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U103 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U104 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U105 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U106 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U107 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U108 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U109 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U110 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U111 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U112 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U113 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U114 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U115 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U116 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U117 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U118 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U119 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U120 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U121 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U122 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U123 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U124 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U125 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U126 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U127 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
endmodule


module BWAdder_57 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U3 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U4 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U5 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U6 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U7 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U8 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U9 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U10 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U11 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U12 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U13 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U14 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U15 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U16 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U17 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U18 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U19 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U20 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U21 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U22 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U23 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U24 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U25 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U26 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U27 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U28 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U29 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U30 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U31 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U32 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U33 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U34 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U35 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U36 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U37 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U38 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U39 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U40 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U41 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U42 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U43 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U44 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U45 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U46 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U47 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U48 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U49 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U50 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U51 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U52 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U53 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U54 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U55 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U56 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U57 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U58 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U59 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U60 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U61 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U62 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U63 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U64 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U65 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U66 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U67 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U68 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U69 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U70 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U71 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U72 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U73 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U74 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U75 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U76 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U77 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U78 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U79 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U80 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U81 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U82 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U83 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U84 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U85 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U86 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U87 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U88 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U89 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U90 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U91 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U92 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U93 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U94 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U95 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U96 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U97 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U98 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U99 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U100 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U101 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U102 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U103 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U104 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U105 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U106 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U107 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U108 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U109 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U110 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U111 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U112 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U113 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U114 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U115 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U116 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U117 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U118 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U119 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U120 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U121 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
  INV_X1 U122 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U123 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U124 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U125 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U126 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U127 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
endmodule


module BWAdder_58 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n190), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n189), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n188), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n187), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n187) );
  XOR2_X1 U134 ( .A(c[62]), .B(n186), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n185), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n184), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n183), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n182), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n181), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n180), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n179), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n178), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n177), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n176), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n175), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n174), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n173), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n172), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n171), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n170), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n169), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n168), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n167), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n166), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n165), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n164), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n163), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n162), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n161), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n160), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n159), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n158), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n157), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n156), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n155), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n154), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n153), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n152), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n151), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n150), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n149), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n148), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n147), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n146), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n145), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n144), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n143), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n142), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n141), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n140), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n139), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n138), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n137), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n136), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n135), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n134), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n133), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n132), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n131), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n130), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n129), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n128), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n190) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n189) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n188) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n183) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n186) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n185) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n184) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n182) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n172) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n181) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n180) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n179) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n178) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n177) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n176) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n175) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n174) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n173) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n171) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n161) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n170) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n169) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n168) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n167) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n166) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n165) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n164) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n163) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n162) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n160) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n150) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n159) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n158) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n157) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n156) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n155) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n154) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n153) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n152) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n151) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n149) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n139) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n148) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n147) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n146) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n145) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n144) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n143) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n142) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n141) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n140) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n138) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n128) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n137) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n136) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n135) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n134) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n133) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n132) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n131) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n130) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n129) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n191) );
  INV_X1 U2 ( .A(n8), .ZN(carry[17]) );
  AOI22_X1 U3 ( .A1(b[16]), .A2(a[16]), .B1(n135), .B2(c[16]), .ZN(n8) );
  INV_X1 U4 ( .A(n13), .ZN(carry[21]) );
  AOI22_X1 U5 ( .A1(b[20]), .A2(a[20]), .B1(n140), .B2(c[20]), .ZN(n13) );
  INV_X1 U6 ( .A(n9), .ZN(carry[18]) );
  AOI22_X1 U7 ( .A1(b[17]), .A2(a[17]), .B1(n136), .B2(c[17]), .ZN(n9) );
  INV_X1 U8 ( .A(n7), .ZN(carry[16]) );
  AOI22_X1 U9 ( .A1(b[15]), .A2(a[15]), .B1(n134), .B2(c[15]), .ZN(n7) );
  INV_X1 U10 ( .A(n6), .ZN(carry[15]) );
  AOI22_X1 U11 ( .A1(b[14]), .A2(a[14]), .B1(n133), .B2(c[14]), .ZN(n6) );
  INV_X1 U12 ( .A(n10), .ZN(carry[19]) );
  AOI22_X1 U13 ( .A1(b[18]), .A2(a[18]), .B1(n137), .B2(c[18]), .ZN(n10) );
  INV_X1 U14 ( .A(n12), .ZN(carry[20]) );
  AOI22_X1 U15 ( .A1(b[19]), .A2(a[19]), .B1(n138), .B2(c[19]), .ZN(n12) );
  INV_X1 U16 ( .A(n14), .ZN(carry[22]) );
  AOI22_X1 U17 ( .A1(b[21]), .A2(a[21]), .B1(n141), .B2(c[21]), .ZN(n14) );
  INV_X1 U18 ( .A(n15), .ZN(carry[23]) );
  AOI22_X1 U19 ( .A1(b[22]), .A2(a[22]), .B1(n142), .B2(c[22]), .ZN(n15) );
  INV_X1 U20 ( .A(n16), .ZN(carry[24]) );
  AOI22_X1 U21 ( .A1(b[23]), .A2(a[23]), .B1(n143), .B2(c[23]), .ZN(n16) );
  INV_X1 U22 ( .A(n17), .ZN(carry[25]) );
  AOI22_X1 U23 ( .A1(b[24]), .A2(a[24]), .B1(n144), .B2(c[24]), .ZN(n17) );
  INV_X1 U24 ( .A(n18), .ZN(carry[26]) );
  AOI22_X1 U25 ( .A1(b[25]), .A2(a[25]), .B1(n145), .B2(c[25]), .ZN(n18) );
  INV_X1 U26 ( .A(n19), .ZN(carry[27]) );
  AOI22_X1 U27 ( .A1(b[26]), .A2(a[26]), .B1(n146), .B2(c[26]), .ZN(n19) );
  INV_X1 U28 ( .A(n29), .ZN(carry[36]) );
  AOI22_X1 U29 ( .A1(b[35]), .A2(a[35]), .B1(n156), .B2(c[35]), .ZN(n29) );
  INV_X1 U30 ( .A(n30), .ZN(carry[37]) );
  AOI22_X1 U31 ( .A1(b[36]), .A2(a[36]), .B1(n157), .B2(c[36]), .ZN(n30) );
  INV_X1 U32 ( .A(n31), .ZN(carry[38]) );
  AOI22_X1 U33 ( .A1(b[37]), .A2(a[37]), .B1(n158), .B2(c[37]), .ZN(n31) );
  INV_X1 U34 ( .A(n32), .ZN(carry[39]) );
  AOI22_X1 U35 ( .A1(b[38]), .A2(a[38]), .B1(n159), .B2(c[38]), .ZN(n32) );
  INV_X1 U36 ( .A(n34), .ZN(carry[40]) );
  AOI22_X1 U37 ( .A1(b[39]), .A2(a[39]), .B1(n160), .B2(c[39]), .ZN(n34) );
  INV_X1 U38 ( .A(n20), .ZN(carry[28]) );
  AOI22_X1 U39 ( .A1(b[27]), .A2(a[27]), .B1(n147), .B2(c[27]), .ZN(n20) );
  INV_X1 U40 ( .A(n21), .ZN(carry[29]) );
  AOI22_X1 U41 ( .A1(b[28]), .A2(a[28]), .B1(n148), .B2(c[28]), .ZN(n21) );
  INV_X1 U42 ( .A(n23), .ZN(carry[30]) );
  AOI22_X1 U43 ( .A1(b[29]), .A2(a[29]), .B1(n149), .B2(c[29]), .ZN(n23) );
  INV_X1 U44 ( .A(n24), .ZN(carry[31]) );
  AOI22_X1 U45 ( .A1(b[30]), .A2(a[30]), .B1(n151), .B2(c[30]), .ZN(n24) );
  INV_X1 U46 ( .A(n25), .ZN(carry[32]) );
  AOI22_X1 U47 ( .A1(b[31]), .A2(a[31]), .B1(n152), .B2(c[31]), .ZN(n25) );
  INV_X1 U48 ( .A(n26), .ZN(carry[33]) );
  AOI22_X1 U49 ( .A1(b[32]), .A2(a[32]), .B1(n153), .B2(c[32]), .ZN(n26) );
  INV_X1 U50 ( .A(n27), .ZN(carry[34]) );
  AOI22_X1 U51 ( .A1(b[33]), .A2(a[33]), .B1(n154), .B2(c[33]), .ZN(n27) );
  INV_X1 U52 ( .A(n28), .ZN(carry[35]) );
  AOI22_X1 U53 ( .A1(b[34]), .A2(a[34]), .B1(n155), .B2(c[34]), .ZN(n28) );
  INV_X1 U54 ( .A(n35), .ZN(carry[41]) );
  AOI22_X1 U55 ( .A1(b[40]), .A2(a[40]), .B1(n162), .B2(c[40]), .ZN(n35) );
  INV_X1 U56 ( .A(n36), .ZN(carry[42]) );
  AOI22_X1 U57 ( .A1(b[41]), .A2(a[41]), .B1(n163), .B2(c[41]), .ZN(n36) );
  INV_X1 U58 ( .A(n37), .ZN(carry[43]) );
  AOI22_X1 U59 ( .A1(b[42]), .A2(a[42]), .B1(n164), .B2(c[42]), .ZN(n37) );
  INV_X1 U60 ( .A(n38), .ZN(carry[44]) );
  AOI22_X1 U61 ( .A1(b[43]), .A2(a[43]), .B1(n165), .B2(c[43]), .ZN(n38) );
  INV_X1 U62 ( .A(n39), .ZN(carry[45]) );
  AOI22_X1 U63 ( .A1(b[44]), .A2(a[44]), .B1(n166), .B2(c[44]), .ZN(n39) );
  INV_X1 U64 ( .A(n40), .ZN(carry[46]) );
  AOI22_X1 U65 ( .A1(b[45]), .A2(a[45]), .B1(n167), .B2(c[45]), .ZN(n40) );
  INV_X1 U66 ( .A(n41), .ZN(carry[47]) );
  AOI22_X1 U67 ( .A1(b[46]), .A2(a[46]), .B1(n168), .B2(c[46]), .ZN(n41) );
  INV_X1 U68 ( .A(n42), .ZN(carry[48]) );
  AOI22_X1 U69 ( .A1(b[47]), .A2(a[47]), .B1(n169), .B2(c[47]), .ZN(n42) );
  INV_X1 U70 ( .A(n43), .ZN(carry[49]) );
  AOI22_X1 U71 ( .A1(b[48]), .A2(a[48]), .B1(n170), .B2(c[48]), .ZN(n43) );
  INV_X1 U72 ( .A(n45), .ZN(carry[50]) );
  AOI22_X1 U73 ( .A1(b[49]), .A2(a[49]), .B1(n171), .B2(c[49]), .ZN(n45) );
  INV_X1 U74 ( .A(n46), .ZN(carry[51]) );
  AOI22_X1 U75 ( .A1(b[50]), .A2(a[50]), .B1(n173), .B2(c[50]), .ZN(n46) );
  INV_X1 U76 ( .A(n47), .ZN(carry[52]) );
  AOI22_X1 U77 ( .A1(b[51]), .A2(a[51]), .B1(n174), .B2(c[51]), .ZN(n47) );
  INV_X1 U78 ( .A(n48), .ZN(carry[53]) );
  AOI22_X1 U79 ( .A1(b[52]), .A2(a[52]), .B1(n175), .B2(c[52]), .ZN(n48) );
  INV_X1 U80 ( .A(n49), .ZN(carry[54]) );
  AOI22_X1 U81 ( .A1(b[53]), .A2(a[53]), .B1(n176), .B2(c[53]), .ZN(n49) );
  INV_X1 U82 ( .A(n52), .ZN(carry[57]) );
  AOI22_X1 U83 ( .A1(b[56]), .A2(a[56]), .B1(n179), .B2(c[56]), .ZN(n52) );
  INV_X1 U84 ( .A(n54), .ZN(carry[59]) );
  AOI22_X1 U85 ( .A1(b[58]), .A2(a[58]), .B1(n181), .B2(c[58]), .ZN(n54) );
  INV_X1 U86 ( .A(n56), .ZN(carry[60]) );
  AOI22_X1 U87 ( .A1(b[59]), .A2(a[59]), .B1(n182), .B2(c[59]), .ZN(n56) );
  INV_X1 U88 ( .A(n57), .ZN(carry[61]) );
  AOI22_X1 U89 ( .A1(b[60]), .A2(a[60]), .B1(n184), .B2(c[60]), .ZN(n57) );
  INV_X1 U90 ( .A(n58), .ZN(carry[62]) );
  AOI22_X1 U91 ( .A1(b[61]), .A2(a[61]), .B1(n185), .B2(c[61]), .ZN(n58) );
  INV_X1 U92 ( .A(n50), .ZN(carry[55]) );
  AOI22_X1 U93 ( .A1(b[54]), .A2(a[54]), .B1(n177), .B2(c[54]), .ZN(n50) );
  INV_X1 U94 ( .A(n51), .ZN(carry[56]) );
  AOI22_X1 U95 ( .A1(b[55]), .A2(a[55]), .B1(n178), .B2(c[55]), .ZN(n51) );
  INV_X1 U96 ( .A(n53), .ZN(carry[58]) );
  AOI22_X1 U97 ( .A1(b[57]), .A2(a[57]), .B1(n180), .B2(c[57]), .ZN(n53) );
  INV_X1 U98 ( .A(n59), .ZN(carry[63]) );
  AOI22_X1 U99 ( .A1(b[62]), .A2(a[62]), .B1(n186), .B2(c[62]), .ZN(n59) );
  INV_X1 U100 ( .A(n5), .ZN(carry[14]) );
  AOI22_X1 U101 ( .A1(b[13]), .A2(a[13]), .B1(n132), .B2(c[13]), .ZN(n5) );
  INV_X1 U102 ( .A(n11), .ZN(carry[1]) );
  AOI22_X1 U103 ( .A1(b[0]), .A2(a[0]), .B1(n128), .B2(c[0]), .ZN(n11) );
  INV_X1 U104 ( .A(n22), .ZN(carry[2]) );
  AOI22_X1 U105 ( .A1(b[1]), .A2(a[1]), .B1(n139), .B2(c[1]), .ZN(n22) );
  INV_X1 U106 ( .A(n33), .ZN(carry[3]) );
  AOI22_X1 U107 ( .A1(b[2]), .A2(a[2]), .B1(n150), .B2(c[2]), .ZN(n33) );
  INV_X1 U108 ( .A(n44), .ZN(carry[4]) );
  AOI22_X1 U109 ( .A1(b[3]), .A2(a[3]), .B1(n161), .B2(c[3]), .ZN(n44) );
  INV_X1 U110 ( .A(n55), .ZN(carry[5]) );
  AOI22_X1 U111 ( .A1(b[4]), .A2(a[4]), .B1(n172), .B2(c[4]), .ZN(n55) );
  INV_X1 U112 ( .A(n60), .ZN(carry[6]) );
  AOI22_X1 U113 ( .A1(b[5]), .A2(a[5]), .B1(n183), .B2(c[5]), .ZN(n60) );
  INV_X1 U114 ( .A(n61), .ZN(carry[7]) );
  AOI22_X1 U115 ( .A1(b[6]), .A2(a[6]), .B1(n188), .B2(c[6]), .ZN(n61) );
  INV_X1 U116 ( .A(n62), .ZN(carry[8]) );
  AOI22_X1 U117 ( .A1(b[7]), .A2(a[7]), .B1(n189), .B2(c[7]), .ZN(n62) );
  INV_X1 U118 ( .A(n63), .ZN(carry[9]) );
  AOI22_X1 U119 ( .A1(b[8]), .A2(a[8]), .B1(n190), .B2(c[8]), .ZN(n63) );
  INV_X1 U120 ( .A(n1), .ZN(carry[10]) );
  AOI22_X1 U121 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n1) );
  INV_X1 U122 ( .A(n2), .ZN(carry[11]) );
  AOI22_X1 U123 ( .A1(b[10]), .A2(a[10]), .B1(n129), .B2(c[10]), .ZN(n2) );
  INV_X1 U124 ( .A(n3), .ZN(carry[12]) );
  AOI22_X1 U125 ( .A1(b[11]), .A2(a[11]), .B1(n130), .B2(c[11]), .ZN(n3) );
  INV_X1 U126 ( .A(n4), .ZN(carry[13]) );
  AOI22_X1 U127 ( .A1(b[12]), .A2(a[12]), .B1(n131), .B2(c[12]), .ZN(n4) );
endmodule


module BWAdder_59 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(c[9]), .B(n193), .Z(result[9]) );
  XOR2_X1 U129 ( .A(c[8]), .B(n192), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n191), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n190), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n189), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n189) );
  XOR2_X1 U134 ( .A(c[62]), .B(n188), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n187), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n186), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n185), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n184), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n183), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n182), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n181), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n180), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n179), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n178), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n177), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n176), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n175), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n174), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n173), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n172), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n171), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n170), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n169), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n168), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n167), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n166), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n165), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n164), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n163), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n162), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n161), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n160), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n159), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n158), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n157), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n156), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n155), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n154), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n153), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n152), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n151), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n150), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n149), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n148), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n147), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n146), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n145), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n144), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n143), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n142), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n141), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n140), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n139), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n138), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n137), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n136), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n135), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n134), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n133), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n132), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n131), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n130), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n192) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n191) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n190) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n185) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n188) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n187) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n186) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n184) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n174) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n183) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n182) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n181) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n180) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n179) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n178) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n177) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n176) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n175) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n173) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n163) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n172) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n171) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n170) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n169) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n168) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n167) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n166) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n165) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n164) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n162) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n152) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n161) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n160) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n159) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n158) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n157) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n156) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n155) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n154) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n153) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n151) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n141) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n150) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n149) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n148) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n147) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n146) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n145) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n144) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n143) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n142) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n140) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n130) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n139) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n138) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n137) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n136) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n135) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n134) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n133) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n132) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n131) );
  INV_X1 U2 ( .A(b[9]), .ZN(n1) );
  XNOR2_X1 U3 ( .A(a[9]), .B(n1), .ZN(n193) );
  INV_X1 U4 ( .A(n14), .ZN(carry[21]) );
  AOI22_X1 U5 ( .A1(b[20]), .A2(a[20]), .B1(n142), .B2(c[20]), .ZN(n14) );
  INV_X1 U6 ( .A(n15), .ZN(carry[22]) );
  AOI22_X1 U7 ( .A1(b[21]), .A2(a[21]), .B1(n143), .B2(c[21]), .ZN(n15) );
  INV_X1 U8 ( .A(n13), .ZN(carry[20]) );
  AOI22_X1 U9 ( .A1(b[19]), .A2(a[19]), .B1(n140), .B2(c[19]), .ZN(n13) );
  INV_X1 U10 ( .A(n7), .ZN(carry[15]) );
  AOI22_X1 U11 ( .A1(b[14]), .A2(a[14]), .B1(n135), .B2(c[14]), .ZN(n7) );
  INV_X1 U12 ( .A(n4), .ZN(carry[12]) );
  AOI22_X1 U13 ( .A1(b[11]), .A2(a[11]), .B1(n132), .B2(c[11]), .ZN(n4) );
  INV_X1 U14 ( .A(n8), .ZN(carry[16]) );
  AOI22_X1 U15 ( .A1(b[15]), .A2(a[15]), .B1(n136), .B2(c[15]), .ZN(n8) );
  INV_X1 U16 ( .A(n9), .ZN(carry[17]) );
  AOI22_X1 U17 ( .A1(b[16]), .A2(a[16]), .B1(n137), .B2(c[16]), .ZN(n9) );
  INV_X1 U18 ( .A(n5), .ZN(carry[13]) );
  AOI22_X1 U19 ( .A1(b[12]), .A2(a[12]), .B1(n133), .B2(c[12]), .ZN(n5) );
  INV_X1 U20 ( .A(n6), .ZN(carry[14]) );
  AOI22_X1 U21 ( .A1(b[13]), .A2(a[13]), .B1(n134), .B2(c[13]), .ZN(n6) );
  INV_X1 U22 ( .A(n10), .ZN(carry[18]) );
  AOI22_X1 U23 ( .A1(b[17]), .A2(a[17]), .B1(n138), .B2(c[17]), .ZN(n10) );
  INV_X1 U24 ( .A(n11), .ZN(carry[19]) );
  AOI22_X1 U25 ( .A1(b[18]), .A2(a[18]), .B1(n139), .B2(c[18]), .ZN(n11) );
  INV_X1 U26 ( .A(n16), .ZN(carry[23]) );
  AOI22_X1 U27 ( .A1(b[22]), .A2(a[22]), .B1(n144), .B2(c[22]), .ZN(n16) );
  INV_X1 U28 ( .A(n17), .ZN(carry[24]) );
  AOI22_X1 U29 ( .A1(b[23]), .A2(a[23]), .B1(n145), .B2(c[23]), .ZN(n17) );
  INV_X1 U30 ( .A(n18), .ZN(carry[25]) );
  AOI22_X1 U31 ( .A1(b[24]), .A2(a[24]), .B1(n146), .B2(c[24]), .ZN(n18) );
  INV_X1 U32 ( .A(n19), .ZN(carry[26]) );
  AOI22_X1 U33 ( .A1(b[25]), .A2(a[25]), .B1(n147), .B2(c[25]), .ZN(n19) );
  INV_X1 U34 ( .A(n20), .ZN(carry[27]) );
  AOI22_X1 U35 ( .A1(b[26]), .A2(a[26]), .B1(n148), .B2(c[26]), .ZN(n20) );
  INV_X1 U36 ( .A(n30), .ZN(carry[36]) );
  AOI22_X1 U37 ( .A1(b[35]), .A2(a[35]), .B1(n158), .B2(c[35]), .ZN(n30) );
  INV_X1 U38 ( .A(n31), .ZN(carry[37]) );
  AOI22_X1 U39 ( .A1(b[36]), .A2(a[36]), .B1(n159), .B2(c[36]), .ZN(n31) );
  INV_X1 U40 ( .A(n32), .ZN(carry[38]) );
  AOI22_X1 U41 ( .A1(b[37]), .A2(a[37]), .B1(n160), .B2(c[37]), .ZN(n32) );
  INV_X1 U42 ( .A(n33), .ZN(carry[39]) );
  AOI22_X1 U43 ( .A1(b[38]), .A2(a[38]), .B1(n161), .B2(c[38]), .ZN(n33) );
  INV_X1 U44 ( .A(n35), .ZN(carry[40]) );
  AOI22_X1 U45 ( .A1(b[39]), .A2(a[39]), .B1(n162), .B2(c[39]), .ZN(n35) );
  INV_X1 U46 ( .A(n21), .ZN(carry[28]) );
  AOI22_X1 U47 ( .A1(b[27]), .A2(a[27]), .B1(n149), .B2(c[27]), .ZN(n21) );
  INV_X1 U48 ( .A(n22), .ZN(carry[29]) );
  AOI22_X1 U49 ( .A1(b[28]), .A2(a[28]), .B1(n150), .B2(c[28]), .ZN(n22) );
  INV_X1 U50 ( .A(n24), .ZN(carry[30]) );
  AOI22_X1 U51 ( .A1(b[29]), .A2(a[29]), .B1(n151), .B2(c[29]), .ZN(n24) );
  INV_X1 U52 ( .A(n25), .ZN(carry[31]) );
  AOI22_X1 U53 ( .A1(b[30]), .A2(a[30]), .B1(n153), .B2(c[30]), .ZN(n25) );
  INV_X1 U54 ( .A(n26), .ZN(carry[32]) );
  AOI22_X1 U55 ( .A1(b[31]), .A2(a[31]), .B1(n154), .B2(c[31]), .ZN(n26) );
  INV_X1 U56 ( .A(n27), .ZN(carry[33]) );
  AOI22_X1 U57 ( .A1(b[32]), .A2(a[32]), .B1(n155), .B2(c[32]), .ZN(n27) );
  INV_X1 U58 ( .A(n28), .ZN(carry[34]) );
  AOI22_X1 U59 ( .A1(b[33]), .A2(a[33]), .B1(n156), .B2(c[33]), .ZN(n28) );
  INV_X1 U60 ( .A(n29), .ZN(carry[35]) );
  AOI22_X1 U61 ( .A1(b[34]), .A2(a[34]), .B1(n157), .B2(c[34]), .ZN(n29) );
  INV_X1 U62 ( .A(n36), .ZN(carry[41]) );
  AOI22_X1 U63 ( .A1(b[40]), .A2(a[40]), .B1(n164), .B2(c[40]), .ZN(n36) );
  INV_X1 U64 ( .A(n37), .ZN(carry[42]) );
  AOI22_X1 U65 ( .A1(b[41]), .A2(a[41]), .B1(n165), .B2(c[41]), .ZN(n37) );
  INV_X1 U66 ( .A(n38), .ZN(carry[43]) );
  AOI22_X1 U67 ( .A1(b[42]), .A2(a[42]), .B1(n166), .B2(c[42]), .ZN(n38) );
  INV_X1 U68 ( .A(n39), .ZN(carry[44]) );
  AOI22_X1 U69 ( .A1(b[43]), .A2(a[43]), .B1(n167), .B2(c[43]), .ZN(n39) );
  INV_X1 U70 ( .A(n40), .ZN(carry[45]) );
  AOI22_X1 U71 ( .A1(b[44]), .A2(a[44]), .B1(n168), .B2(c[44]), .ZN(n40) );
  INV_X1 U72 ( .A(n41), .ZN(carry[46]) );
  AOI22_X1 U73 ( .A1(b[45]), .A2(a[45]), .B1(n169), .B2(c[45]), .ZN(n41) );
  INV_X1 U74 ( .A(n42), .ZN(carry[47]) );
  AOI22_X1 U75 ( .A1(b[46]), .A2(a[46]), .B1(n170), .B2(c[46]), .ZN(n42) );
  INV_X1 U76 ( .A(n43), .ZN(carry[48]) );
  AOI22_X1 U77 ( .A1(b[47]), .A2(a[47]), .B1(n171), .B2(c[47]), .ZN(n43) );
  INV_X1 U78 ( .A(n44), .ZN(carry[49]) );
  AOI22_X1 U79 ( .A1(b[48]), .A2(a[48]), .B1(n172), .B2(c[48]), .ZN(n44) );
  INV_X1 U80 ( .A(n46), .ZN(carry[50]) );
  AOI22_X1 U81 ( .A1(b[49]), .A2(a[49]), .B1(n173), .B2(c[49]), .ZN(n46) );
  INV_X1 U82 ( .A(n47), .ZN(carry[51]) );
  AOI22_X1 U83 ( .A1(b[50]), .A2(a[50]), .B1(n175), .B2(c[50]), .ZN(n47) );
  INV_X1 U84 ( .A(n48), .ZN(carry[52]) );
  AOI22_X1 U85 ( .A1(b[51]), .A2(a[51]), .B1(n176), .B2(c[51]), .ZN(n48) );
  INV_X1 U86 ( .A(n49), .ZN(carry[53]) );
  AOI22_X1 U87 ( .A1(b[52]), .A2(a[52]), .B1(n177), .B2(c[52]), .ZN(n49) );
  INV_X1 U88 ( .A(n50), .ZN(carry[54]) );
  AOI22_X1 U89 ( .A1(b[53]), .A2(a[53]), .B1(n178), .B2(c[53]), .ZN(n50) );
  INV_X1 U90 ( .A(n51), .ZN(carry[55]) );
  AOI22_X1 U91 ( .A1(b[54]), .A2(a[54]), .B1(n179), .B2(c[54]), .ZN(n51) );
  INV_X1 U92 ( .A(n52), .ZN(carry[56]) );
  AOI22_X1 U93 ( .A1(b[55]), .A2(a[55]), .B1(n180), .B2(c[55]), .ZN(n52) );
  INV_X1 U94 ( .A(n53), .ZN(carry[57]) );
  AOI22_X1 U95 ( .A1(b[56]), .A2(a[56]), .B1(n181), .B2(c[56]), .ZN(n53) );
  INV_X1 U96 ( .A(n54), .ZN(carry[58]) );
  AOI22_X1 U97 ( .A1(b[57]), .A2(a[57]), .B1(n182), .B2(c[57]), .ZN(n54) );
  INV_X1 U98 ( .A(n55), .ZN(carry[59]) );
  AOI22_X1 U99 ( .A1(b[58]), .A2(a[58]), .B1(n183), .B2(c[58]), .ZN(n55) );
  INV_X1 U100 ( .A(n57), .ZN(carry[60]) );
  AOI22_X1 U101 ( .A1(b[59]), .A2(a[59]), .B1(n184), .B2(c[59]), .ZN(n57) );
  INV_X1 U102 ( .A(n58), .ZN(carry[61]) );
  AOI22_X1 U103 ( .A1(b[60]), .A2(a[60]), .B1(n186), .B2(c[60]), .ZN(n58) );
  INV_X1 U104 ( .A(n59), .ZN(carry[62]) );
  AOI22_X1 U105 ( .A1(b[61]), .A2(a[61]), .B1(n187), .B2(c[61]), .ZN(n59) );
  INV_X1 U106 ( .A(n60), .ZN(carry[63]) );
  AOI22_X1 U107 ( .A1(b[62]), .A2(a[62]), .B1(n188), .B2(c[62]), .ZN(n60) );
  INV_X1 U108 ( .A(n3), .ZN(carry[11]) );
  INV_X1 U109 ( .A(n12), .ZN(carry[1]) );
  AOI22_X1 U110 ( .A1(b[0]), .A2(a[0]), .B1(n130), .B2(c[0]), .ZN(n12) );
  INV_X1 U111 ( .A(n23), .ZN(carry[2]) );
  AOI22_X1 U112 ( .A1(b[1]), .A2(a[1]), .B1(n141), .B2(c[1]), .ZN(n23) );
  INV_X1 U113 ( .A(n34), .ZN(carry[3]) );
  AOI22_X1 U114 ( .A1(b[2]), .A2(a[2]), .B1(n152), .B2(c[2]), .ZN(n34) );
  INV_X1 U115 ( .A(n45), .ZN(carry[4]) );
  AOI22_X1 U116 ( .A1(b[3]), .A2(a[3]), .B1(n163), .B2(c[3]), .ZN(n45) );
  INV_X1 U117 ( .A(n56), .ZN(carry[5]) );
  AOI22_X1 U118 ( .A1(b[4]), .A2(a[4]), .B1(n174), .B2(c[4]), .ZN(n56) );
  INV_X1 U119 ( .A(n61), .ZN(carry[6]) );
  AOI22_X1 U120 ( .A1(b[5]), .A2(a[5]), .B1(n185), .B2(c[5]), .ZN(n61) );
  INV_X1 U121 ( .A(n62), .ZN(carry[7]) );
  AOI22_X1 U122 ( .A1(b[6]), .A2(a[6]), .B1(n190), .B2(c[6]), .ZN(n62) );
  INV_X1 U123 ( .A(n63), .ZN(carry[8]) );
  AOI22_X1 U124 ( .A1(b[7]), .A2(a[7]), .B1(n191), .B2(c[7]), .ZN(n63) );
  INV_X1 U125 ( .A(n129), .ZN(carry[9]) );
  AOI22_X1 U126 ( .A1(b[8]), .A2(a[8]), .B1(n192), .B2(c[8]), .ZN(n129) );
  INV_X1 U127 ( .A(n2), .ZN(carry[10]) );
  AOI22_X1 U255 ( .A1(b[9]), .A2(a[9]), .B1(n193), .B2(c[9]), .ZN(n2) );
  AOI22_X1 U256 ( .A1(b[10]), .A2(a[10]), .B1(n131), .B2(c[10]), .ZN(n3) );
endmodule


module BWAdder_60 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(n193), .B(c[9]), .Z(result[9]) );
  XOR2_X1 U129 ( .A(n192), .B(c[8]), .Z(result[8]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n191), .Z(result[7]) );
  XOR2_X1 U131 ( .A(c[6]), .B(n190), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n189), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n189) );
  XOR2_X1 U134 ( .A(c[62]), .B(n188), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n187), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n186), .Z(result[60]) );
  XOR2_X1 U137 ( .A(c[5]), .B(n185), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n184), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n183), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n182), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n181), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n180), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n179), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n178), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n177), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n176), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n175), .Z(result[50]) );
  XOR2_X1 U148 ( .A(c[4]), .B(n174), .Z(result[4]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n173), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n172), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n171), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n170), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n169), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n168), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n167), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n166), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n165), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n164), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n163), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n162), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n161), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n160), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n159), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n158), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n157), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n156), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n155), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n154), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n153), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n152), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n151), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n150), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n149), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n148), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n147), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n146), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n145), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n144), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n143), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n142), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n141), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n140), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n139), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n138), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n137), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n136), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n135), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n134), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n133), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n132), .Z(result[11]) );
  XOR2_X1 U191 ( .A(c[10]), .B(n131), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n130), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n192) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n191) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n190) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n185) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n188) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n187) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n186) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n184) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n174) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n183) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n182) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n181) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n180) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n179) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n178) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n177) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n176) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n175) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n173) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n163) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n172) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n171) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n170) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n169) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n168) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n167) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n166) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n165) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n164) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n162) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n152) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n161) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n160) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n159) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n158) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n157) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n156) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n155) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n154) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n153) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n151) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n141) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n150) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n149) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n148) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n147) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n146) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n145) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n144) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n143) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n142) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n140) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n130) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n139) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n138) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n137) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n136) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n135) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n134) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n133) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n132) );
  XOR2_X1 U254 ( .A(a[10]), .B(b[10]), .Z(n131) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n193) );
  CLKBUF_X1 U2 ( .A(a[8]), .Z(n1) );
  INV_X1 U3 ( .A(n8), .ZN(carry[16]) );
  AOI22_X1 U4 ( .A1(b[15]), .A2(a[15]), .B1(n136), .B2(c[15]), .ZN(n8) );
  INV_X1 U5 ( .A(n129), .ZN(carry[9]) );
  AOI22_X1 U6 ( .A1(b[8]), .A2(n1), .B1(n192), .B2(c[8]), .ZN(n129) );
  INV_X1 U7 ( .A(n2), .ZN(carry[10]) );
  AOI22_X1 U8 ( .A1(b[9]), .A2(a[9]), .B1(n193), .B2(c[9]), .ZN(n2) );
  INV_X1 U9 ( .A(n9), .ZN(carry[17]) );
  AOI22_X1 U10 ( .A1(b[16]), .A2(a[16]), .B1(n137), .B2(c[16]), .ZN(n9) );
  INV_X1 U11 ( .A(n3), .ZN(carry[11]) );
  AOI22_X1 U12 ( .A1(b[10]), .A2(a[10]), .B1(n131), .B2(c[10]), .ZN(n3) );
  INV_X1 U13 ( .A(n4), .ZN(carry[12]) );
  AOI22_X1 U14 ( .A1(b[11]), .A2(a[11]), .B1(n132), .B2(c[11]), .ZN(n4) );
  INV_X1 U15 ( .A(n5), .ZN(carry[13]) );
  AOI22_X1 U16 ( .A1(b[12]), .A2(a[12]), .B1(n133), .B2(c[12]), .ZN(n5) );
  INV_X1 U17 ( .A(n6), .ZN(carry[14]) );
  AOI22_X1 U18 ( .A1(b[13]), .A2(a[13]), .B1(n134), .B2(c[13]), .ZN(n6) );
  INV_X1 U19 ( .A(n7), .ZN(carry[15]) );
  AOI22_X1 U20 ( .A1(b[14]), .A2(a[14]), .B1(n135), .B2(c[14]), .ZN(n7) );
  INV_X1 U21 ( .A(n10), .ZN(carry[18]) );
  AOI22_X1 U22 ( .A1(b[17]), .A2(a[17]), .B1(n138), .B2(c[17]), .ZN(n10) );
  INV_X1 U23 ( .A(n11), .ZN(carry[19]) );
  AOI22_X1 U24 ( .A1(b[18]), .A2(a[18]), .B1(n139), .B2(c[18]), .ZN(n11) );
  INV_X1 U25 ( .A(n13), .ZN(carry[20]) );
  AOI22_X1 U26 ( .A1(b[19]), .A2(a[19]), .B1(n140), .B2(c[19]), .ZN(n13) );
  INV_X1 U27 ( .A(n14), .ZN(carry[21]) );
  AOI22_X1 U28 ( .A1(b[20]), .A2(a[20]), .B1(n142), .B2(c[20]), .ZN(n14) );
  INV_X1 U29 ( .A(n15), .ZN(carry[22]) );
  AOI22_X1 U30 ( .A1(b[21]), .A2(a[21]), .B1(n143), .B2(c[21]), .ZN(n15) );
  INV_X1 U31 ( .A(n16), .ZN(carry[23]) );
  AOI22_X1 U32 ( .A1(b[22]), .A2(a[22]), .B1(n144), .B2(c[22]), .ZN(n16) );
  INV_X1 U33 ( .A(n17), .ZN(carry[24]) );
  AOI22_X1 U34 ( .A1(b[23]), .A2(a[23]), .B1(n145), .B2(c[23]), .ZN(n17) );
  INV_X1 U35 ( .A(n18), .ZN(carry[25]) );
  AOI22_X1 U36 ( .A1(b[24]), .A2(a[24]), .B1(n146), .B2(c[24]), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(carry[26]) );
  AOI22_X1 U38 ( .A1(b[25]), .A2(a[25]), .B1(n147), .B2(c[25]), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(carry[27]) );
  AOI22_X1 U40 ( .A1(b[26]), .A2(a[26]), .B1(n148), .B2(c[26]), .ZN(n20) );
  INV_X1 U41 ( .A(n26), .ZN(carry[32]) );
  AOI22_X1 U42 ( .A1(b[31]), .A2(a[31]), .B1(n154), .B2(c[31]), .ZN(n26) );
  INV_X1 U43 ( .A(n27), .ZN(carry[33]) );
  AOI22_X1 U44 ( .A1(b[32]), .A2(a[32]), .B1(n155), .B2(c[32]), .ZN(n27) );
  INV_X1 U45 ( .A(n28), .ZN(carry[34]) );
  AOI22_X1 U46 ( .A1(b[33]), .A2(a[33]), .B1(n156), .B2(c[33]), .ZN(n28) );
  INV_X1 U47 ( .A(n30), .ZN(carry[36]) );
  AOI22_X1 U48 ( .A1(b[35]), .A2(a[35]), .B1(n158), .B2(c[35]), .ZN(n30) );
  INV_X1 U49 ( .A(n31), .ZN(carry[37]) );
  AOI22_X1 U50 ( .A1(b[36]), .A2(a[36]), .B1(n159), .B2(c[36]), .ZN(n31) );
  INV_X1 U51 ( .A(n21), .ZN(carry[28]) );
  AOI22_X1 U52 ( .A1(b[27]), .A2(a[27]), .B1(n149), .B2(c[27]), .ZN(n21) );
  INV_X1 U53 ( .A(n22), .ZN(carry[29]) );
  AOI22_X1 U54 ( .A1(b[28]), .A2(a[28]), .B1(n150), .B2(c[28]), .ZN(n22) );
  INV_X1 U55 ( .A(n24), .ZN(carry[30]) );
  AOI22_X1 U56 ( .A1(b[29]), .A2(a[29]), .B1(n151), .B2(c[29]), .ZN(n24) );
  INV_X1 U57 ( .A(n25), .ZN(carry[31]) );
  AOI22_X1 U58 ( .A1(b[30]), .A2(a[30]), .B1(n153), .B2(c[30]), .ZN(n25) );
  INV_X1 U59 ( .A(n29), .ZN(carry[35]) );
  AOI22_X1 U60 ( .A1(b[34]), .A2(a[34]), .B1(n157), .B2(c[34]), .ZN(n29) );
  INV_X1 U61 ( .A(n32), .ZN(carry[38]) );
  AOI22_X1 U62 ( .A1(b[37]), .A2(a[37]), .B1(n160), .B2(c[37]), .ZN(n32) );
  INV_X1 U63 ( .A(n33), .ZN(carry[39]) );
  AOI22_X1 U64 ( .A1(b[38]), .A2(a[38]), .B1(n161), .B2(c[38]), .ZN(n33) );
  INV_X1 U65 ( .A(n35), .ZN(carry[40]) );
  AOI22_X1 U66 ( .A1(b[39]), .A2(a[39]), .B1(n162), .B2(c[39]), .ZN(n35) );
  INV_X1 U67 ( .A(n36), .ZN(carry[41]) );
  AOI22_X1 U68 ( .A1(b[40]), .A2(a[40]), .B1(n164), .B2(c[40]), .ZN(n36) );
  INV_X1 U69 ( .A(n37), .ZN(carry[42]) );
  AOI22_X1 U70 ( .A1(b[41]), .A2(a[41]), .B1(n165), .B2(c[41]), .ZN(n37) );
  INV_X1 U71 ( .A(n38), .ZN(carry[43]) );
  AOI22_X1 U72 ( .A1(b[42]), .A2(a[42]), .B1(n166), .B2(c[42]), .ZN(n38) );
  INV_X1 U73 ( .A(n39), .ZN(carry[44]) );
  AOI22_X1 U74 ( .A1(b[43]), .A2(a[43]), .B1(n167), .B2(c[43]), .ZN(n39) );
  INV_X1 U75 ( .A(n40), .ZN(carry[45]) );
  AOI22_X1 U76 ( .A1(b[44]), .A2(a[44]), .B1(n168), .B2(c[44]), .ZN(n40) );
  INV_X1 U77 ( .A(n41), .ZN(carry[46]) );
  AOI22_X1 U78 ( .A1(b[45]), .A2(a[45]), .B1(n169), .B2(c[45]), .ZN(n41) );
  INV_X1 U79 ( .A(n42), .ZN(carry[47]) );
  AOI22_X1 U80 ( .A1(b[46]), .A2(a[46]), .B1(n170), .B2(c[46]), .ZN(n42) );
  INV_X1 U81 ( .A(n43), .ZN(carry[48]) );
  AOI22_X1 U82 ( .A1(b[47]), .A2(a[47]), .B1(n171), .B2(c[47]), .ZN(n43) );
  INV_X1 U83 ( .A(n44), .ZN(carry[49]) );
  AOI22_X1 U84 ( .A1(b[48]), .A2(a[48]), .B1(n172), .B2(c[48]), .ZN(n44) );
  INV_X1 U85 ( .A(n46), .ZN(carry[50]) );
  AOI22_X1 U86 ( .A1(b[49]), .A2(a[49]), .B1(n173), .B2(c[49]), .ZN(n46) );
  INV_X1 U87 ( .A(n47), .ZN(carry[51]) );
  AOI22_X1 U88 ( .A1(b[50]), .A2(a[50]), .B1(n175), .B2(c[50]), .ZN(n47) );
  INV_X1 U89 ( .A(n48), .ZN(carry[52]) );
  AOI22_X1 U90 ( .A1(b[51]), .A2(a[51]), .B1(n176), .B2(c[51]), .ZN(n48) );
  INV_X1 U91 ( .A(n49), .ZN(carry[53]) );
  AOI22_X1 U92 ( .A1(b[52]), .A2(a[52]), .B1(n177), .B2(c[52]), .ZN(n49) );
  INV_X1 U93 ( .A(n50), .ZN(carry[54]) );
  AOI22_X1 U94 ( .A1(b[53]), .A2(a[53]), .B1(n178), .B2(c[53]), .ZN(n50) );
  INV_X1 U95 ( .A(n51), .ZN(carry[55]) );
  AOI22_X1 U96 ( .A1(b[54]), .A2(a[54]), .B1(n179), .B2(c[54]), .ZN(n51) );
  INV_X1 U97 ( .A(n52), .ZN(carry[56]) );
  AOI22_X1 U98 ( .A1(b[55]), .A2(a[55]), .B1(n180), .B2(c[55]), .ZN(n52) );
  INV_X1 U99 ( .A(n53), .ZN(carry[57]) );
  AOI22_X1 U100 ( .A1(b[56]), .A2(a[56]), .B1(n181), .B2(c[56]), .ZN(n53) );
  INV_X1 U101 ( .A(n54), .ZN(carry[58]) );
  AOI22_X1 U102 ( .A1(b[57]), .A2(a[57]), .B1(n182), .B2(c[57]), .ZN(n54) );
  INV_X1 U103 ( .A(n55), .ZN(carry[59]) );
  AOI22_X1 U104 ( .A1(b[58]), .A2(a[58]), .B1(n183), .B2(c[58]), .ZN(n55) );
  INV_X1 U105 ( .A(n57), .ZN(carry[60]) );
  AOI22_X1 U106 ( .A1(b[59]), .A2(a[59]), .B1(n184), .B2(c[59]), .ZN(n57) );
  INV_X1 U107 ( .A(n58), .ZN(carry[61]) );
  AOI22_X1 U108 ( .A1(b[60]), .A2(a[60]), .B1(n186), .B2(c[60]), .ZN(n58) );
  INV_X1 U109 ( .A(n59), .ZN(carry[62]) );
  AOI22_X1 U110 ( .A1(b[61]), .A2(a[61]), .B1(n187), .B2(c[61]), .ZN(n59) );
  INV_X1 U111 ( .A(n60), .ZN(carry[63]) );
  AOI22_X1 U112 ( .A1(b[62]), .A2(a[62]), .B1(n188), .B2(c[62]), .ZN(n60) );
  INV_X1 U113 ( .A(n63), .ZN(carry[8]) );
  AOI22_X1 U114 ( .A1(b[7]), .A2(a[7]), .B1(n191), .B2(c[7]), .ZN(n63) );
  INV_X1 U115 ( .A(n12), .ZN(carry[1]) );
  AOI22_X1 U116 ( .A1(b[0]), .A2(a[0]), .B1(n130), .B2(c[0]), .ZN(n12) );
  INV_X1 U117 ( .A(n23), .ZN(carry[2]) );
  AOI22_X1 U118 ( .A1(b[1]), .A2(a[1]), .B1(n141), .B2(c[1]), .ZN(n23) );
  INV_X1 U119 ( .A(n34), .ZN(carry[3]) );
  AOI22_X1 U120 ( .A1(b[2]), .A2(a[2]), .B1(n152), .B2(c[2]), .ZN(n34) );
  INV_X1 U121 ( .A(n45), .ZN(carry[4]) );
  AOI22_X1 U122 ( .A1(b[3]), .A2(a[3]), .B1(n163), .B2(c[3]), .ZN(n45) );
  INV_X1 U123 ( .A(n56), .ZN(carry[5]) );
  AOI22_X1 U124 ( .A1(b[4]), .A2(a[4]), .B1(n174), .B2(c[4]), .ZN(n56) );
  INV_X1 U125 ( .A(n61), .ZN(carry[6]) );
  AOI22_X1 U126 ( .A1(b[5]), .A2(a[5]), .B1(n185), .B2(c[5]), .ZN(n61) );
  INV_X1 U127 ( .A(n62), .ZN(carry[7]) );
  AOI22_X1 U256 ( .A1(b[6]), .A2(a[6]), .B1(n190), .B2(c[6]), .ZN(n62) );
endmodule


module BWAdder_61 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213;
  assign carry[0] = 1'b0;

  XOR2_X1 U128 ( .A(n213), .B(c[9]), .Z(result[9]) );
  XOR2_X1 U130 ( .A(c[7]), .B(n211), .Z(result[7]) );
  XOR2_X1 U131 ( .A(n210), .B(c[6]), .Z(result[6]) );
  XOR2_X1 U132 ( .A(a[63]), .B(n209), .Z(result[63]) );
  XOR2_X1 U133 ( .A(c[63]), .B(b[63]), .Z(n209) );
  XOR2_X1 U134 ( .A(c[62]), .B(n208), .Z(result[62]) );
  XOR2_X1 U135 ( .A(c[61]), .B(n207), .Z(result[61]) );
  XOR2_X1 U136 ( .A(c[60]), .B(n206), .Z(result[60]) );
  XOR2_X1 U137 ( .A(n205), .B(c[5]), .Z(result[5]) );
  XOR2_X1 U138 ( .A(c[59]), .B(n204), .Z(result[59]) );
  XOR2_X1 U139 ( .A(c[58]), .B(n203), .Z(result[58]) );
  XOR2_X1 U140 ( .A(c[57]), .B(n202), .Z(result[57]) );
  XOR2_X1 U141 ( .A(c[56]), .B(n201), .Z(result[56]) );
  XOR2_X1 U142 ( .A(c[55]), .B(n200), .Z(result[55]) );
  XOR2_X1 U143 ( .A(c[54]), .B(n199), .Z(result[54]) );
  XOR2_X1 U144 ( .A(c[53]), .B(n198), .Z(result[53]) );
  XOR2_X1 U145 ( .A(c[52]), .B(n197), .Z(result[52]) );
  XOR2_X1 U146 ( .A(c[51]), .B(n196), .Z(result[51]) );
  XOR2_X1 U147 ( .A(c[50]), .B(n195), .Z(result[50]) );
  XOR2_X1 U149 ( .A(c[49]), .B(n193), .Z(result[49]) );
  XOR2_X1 U150 ( .A(c[48]), .B(n192), .Z(result[48]) );
  XOR2_X1 U151 ( .A(c[47]), .B(n191), .Z(result[47]) );
  XOR2_X1 U152 ( .A(c[46]), .B(n190), .Z(result[46]) );
  XOR2_X1 U153 ( .A(c[45]), .B(n189), .Z(result[45]) );
  XOR2_X1 U154 ( .A(c[44]), .B(n188), .Z(result[44]) );
  XOR2_X1 U155 ( .A(c[43]), .B(n187), .Z(result[43]) );
  XOR2_X1 U156 ( .A(c[42]), .B(n186), .Z(result[42]) );
  XOR2_X1 U157 ( .A(c[41]), .B(n185), .Z(result[41]) );
  XOR2_X1 U158 ( .A(c[40]), .B(n184), .Z(result[40]) );
  XOR2_X1 U159 ( .A(c[3]), .B(n183), .Z(result[3]) );
  XOR2_X1 U160 ( .A(c[39]), .B(n182), .Z(result[39]) );
  XOR2_X1 U161 ( .A(c[38]), .B(n181), .Z(result[38]) );
  XOR2_X1 U162 ( .A(c[37]), .B(n180), .Z(result[37]) );
  XOR2_X1 U163 ( .A(c[36]), .B(n179), .Z(result[36]) );
  XOR2_X1 U164 ( .A(c[35]), .B(n178), .Z(result[35]) );
  XOR2_X1 U165 ( .A(c[34]), .B(n177), .Z(result[34]) );
  XOR2_X1 U166 ( .A(c[33]), .B(n176), .Z(result[33]) );
  XOR2_X1 U167 ( .A(c[32]), .B(n175), .Z(result[32]) );
  XOR2_X1 U168 ( .A(c[31]), .B(n174), .Z(result[31]) );
  XOR2_X1 U169 ( .A(c[30]), .B(n173), .Z(result[30]) );
  XOR2_X1 U170 ( .A(c[2]), .B(n172), .Z(result[2]) );
  XOR2_X1 U171 ( .A(c[29]), .B(n171), .Z(result[29]) );
  XOR2_X1 U172 ( .A(c[28]), .B(n170), .Z(result[28]) );
  XOR2_X1 U173 ( .A(c[27]), .B(n169), .Z(result[27]) );
  XOR2_X1 U174 ( .A(c[26]), .B(n168), .Z(result[26]) );
  XOR2_X1 U175 ( .A(c[25]), .B(n167), .Z(result[25]) );
  XOR2_X1 U176 ( .A(c[24]), .B(n166), .Z(result[24]) );
  XOR2_X1 U177 ( .A(c[23]), .B(n165), .Z(result[23]) );
  XOR2_X1 U178 ( .A(c[22]), .B(n164), .Z(result[22]) );
  XOR2_X1 U179 ( .A(c[21]), .B(n163), .Z(result[21]) );
  XOR2_X1 U180 ( .A(c[20]), .B(n162), .Z(result[20]) );
  XOR2_X1 U181 ( .A(c[1]), .B(n161), .Z(result[1]) );
  XOR2_X1 U182 ( .A(c[19]), .B(n160), .Z(result[19]) );
  XOR2_X1 U183 ( .A(c[18]), .B(n159), .Z(result[18]) );
  XOR2_X1 U184 ( .A(c[17]), .B(n158), .Z(result[17]) );
  XOR2_X1 U185 ( .A(c[16]), .B(n157), .Z(result[16]) );
  XOR2_X1 U186 ( .A(c[15]), .B(n156), .Z(result[15]) );
  XOR2_X1 U187 ( .A(c[14]), .B(n155), .Z(result[14]) );
  XOR2_X1 U188 ( .A(c[13]), .B(n154), .Z(result[13]) );
  XOR2_X1 U189 ( .A(c[12]), .B(n153), .Z(result[12]) );
  XOR2_X1 U190 ( .A(c[11]), .B(n152), .Z(result[11]) );
  XOR2_X1 U191 ( .A(n151), .B(c[10]), .Z(result[10]) );
  XOR2_X1 U192 ( .A(c[0]), .B(n150), .Z(result[0]) );
  XOR2_X1 U193 ( .A(a[8]), .B(b[8]), .Z(n212) );
  XOR2_X1 U194 ( .A(a[7]), .B(b[7]), .Z(n211) );
  XOR2_X1 U195 ( .A(a[6]), .B(b[6]), .Z(n210) );
  XOR2_X1 U196 ( .A(a[5]), .B(b[5]), .Z(n205) );
  XOR2_X1 U197 ( .A(a[62]), .B(b[62]), .Z(n208) );
  XOR2_X1 U198 ( .A(a[61]), .B(b[61]), .Z(n207) );
  XOR2_X1 U199 ( .A(a[60]), .B(b[60]), .Z(n206) );
  XOR2_X1 U200 ( .A(a[59]), .B(b[59]), .Z(n204) );
  XOR2_X1 U201 ( .A(a[4]), .B(b[4]), .Z(n194) );
  XOR2_X1 U202 ( .A(a[58]), .B(b[58]), .Z(n203) );
  XOR2_X1 U203 ( .A(a[57]), .B(b[57]), .Z(n202) );
  XOR2_X1 U204 ( .A(a[56]), .B(b[56]), .Z(n201) );
  XOR2_X1 U205 ( .A(a[55]), .B(b[55]), .Z(n200) );
  XOR2_X1 U206 ( .A(a[54]), .B(b[54]), .Z(n199) );
  XOR2_X1 U207 ( .A(a[53]), .B(b[53]), .Z(n198) );
  XOR2_X1 U208 ( .A(a[52]), .B(b[52]), .Z(n197) );
  XOR2_X1 U209 ( .A(a[51]), .B(b[51]), .Z(n196) );
  XOR2_X1 U210 ( .A(a[50]), .B(b[50]), .Z(n195) );
  XOR2_X1 U211 ( .A(a[49]), .B(b[49]), .Z(n193) );
  XOR2_X1 U212 ( .A(a[3]), .B(b[3]), .Z(n183) );
  XOR2_X1 U213 ( .A(a[48]), .B(b[48]), .Z(n192) );
  XOR2_X1 U214 ( .A(a[47]), .B(b[47]), .Z(n191) );
  XOR2_X1 U215 ( .A(a[46]), .B(b[46]), .Z(n190) );
  XOR2_X1 U216 ( .A(a[45]), .B(b[45]), .Z(n189) );
  XOR2_X1 U217 ( .A(a[44]), .B(b[44]), .Z(n188) );
  XOR2_X1 U218 ( .A(a[43]), .B(b[43]), .Z(n187) );
  XOR2_X1 U219 ( .A(a[42]), .B(b[42]), .Z(n186) );
  XOR2_X1 U220 ( .A(a[41]), .B(b[41]), .Z(n185) );
  XOR2_X1 U221 ( .A(a[40]), .B(b[40]), .Z(n184) );
  XOR2_X1 U222 ( .A(a[39]), .B(b[39]), .Z(n182) );
  XOR2_X1 U223 ( .A(a[2]), .B(b[2]), .Z(n172) );
  XOR2_X1 U224 ( .A(a[38]), .B(b[38]), .Z(n181) );
  XOR2_X1 U225 ( .A(a[37]), .B(b[37]), .Z(n180) );
  XOR2_X1 U226 ( .A(a[36]), .B(b[36]), .Z(n179) );
  XOR2_X1 U227 ( .A(a[35]), .B(b[35]), .Z(n178) );
  XOR2_X1 U228 ( .A(a[34]), .B(b[34]), .Z(n177) );
  XOR2_X1 U229 ( .A(a[33]), .B(b[33]), .Z(n176) );
  XOR2_X1 U230 ( .A(a[32]), .B(b[32]), .Z(n175) );
  XOR2_X1 U231 ( .A(a[31]), .B(b[31]), .Z(n174) );
  XOR2_X1 U232 ( .A(a[30]), .B(b[30]), .Z(n173) );
  XOR2_X1 U233 ( .A(a[29]), .B(b[29]), .Z(n171) );
  XOR2_X1 U234 ( .A(a[1]), .B(b[1]), .Z(n161) );
  XOR2_X1 U235 ( .A(a[28]), .B(b[28]), .Z(n170) );
  XOR2_X1 U236 ( .A(a[27]), .B(b[27]), .Z(n169) );
  XOR2_X1 U237 ( .A(a[26]), .B(b[26]), .Z(n168) );
  XOR2_X1 U238 ( .A(a[25]), .B(b[25]), .Z(n167) );
  XOR2_X1 U239 ( .A(a[24]), .B(b[24]), .Z(n166) );
  XOR2_X1 U240 ( .A(a[23]), .B(b[23]), .Z(n165) );
  XOR2_X1 U241 ( .A(a[22]), .B(b[22]), .Z(n164) );
  XOR2_X1 U242 ( .A(a[21]), .B(b[21]), .Z(n163) );
  XOR2_X1 U243 ( .A(a[20]), .B(b[20]), .Z(n162) );
  XOR2_X1 U244 ( .A(a[19]), .B(b[19]), .Z(n160) );
  XOR2_X1 U245 ( .A(a[0]), .B(b[0]), .Z(n150) );
  XOR2_X1 U246 ( .A(a[18]), .B(b[18]), .Z(n159) );
  XOR2_X1 U247 ( .A(a[17]), .B(b[17]), .Z(n158) );
  XOR2_X1 U248 ( .A(a[16]), .B(b[16]), .Z(n157) );
  XOR2_X1 U249 ( .A(a[15]), .B(b[15]), .Z(n156) );
  XOR2_X1 U250 ( .A(a[14]), .B(b[14]), .Z(n155) );
  XOR2_X1 U251 ( .A(a[13]), .B(b[13]), .Z(n154) );
  XOR2_X1 U252 ( .A(a[12]), .B(b[12]), .Z(n153) );
  XOR2_X1 U253 ( .A(a[11]), .B(b[11]), .Z(n152) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n213) );
  INV_X1 U2 ( .A(c[4]), .ZN(n6) );
  NAND2_X1 U3 ( .A1(a[10]), .A2(n2), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n1), .A2(b[10]), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n3), .A2(n4), .ZN(n151) );
  INV_X1 U6 ( .A(a[10]), .ZN(n1) );
  INV_X1 U7 ( .A(b[10]), .ZN(n2) );
  CLKBUF_X1 U8 ( .A(a[5]), .Z(n5) );
  XNOR2_X1 U9 ( .A(n194), .B(n6), .ZN(result[4]) );
  INV_X1 U10 ( .A(n23), .ZN(carry[20]) );
  AOI22_X1 U11 ( .A1(b[19]), .A2(a[19]), .B1(n160), .B2(c[19]), .ZN(n23) );
  INV_X1 U12 ( .A(n21), .ZN(carry[19]) );
  AOI22_X1 U13 ( .A1(b[18]), .A2(a[18]), .B1(n159), .B2(c[18]), .ZN(n21) );
  INV_X1 U14 ( .A(n24), .ZN(carry[21]) );
  AOI22_X1 U15 ( .A1(b[20]), .A2(a[20]), .B1(n162), .B2(c[20]), .ZN(n24) );
  INV_X1 U16 ( .A(n30), .ZN(carry[27]) );
  AOI22_X1 U17 ( .A1(b[26]), .A2(a[26]), .B1(n168), .B2(c[26]), .ZN(n30) );
  INV_X1 U18 ( .A(n32), .ZN(carry[29]) );
  AOI22_X1 U19 ( .A1(b[28]), .A2(a[28]), .B1(n170), .B2(c[28]), .ZN(n32) );
  INV_X1 U20 ( .A(n19), .ZN(carry[17]) );
  AOI22_X1 U21 ( .A1(b[16]), .A2(a[16]), .B1(n157), .B2(c[16]), .ZN(n19) );
  INV_X1 U22 ( .A(n13), .ZN(carry[11]) );
  AOI22_X1 U23 ( .A1(b[10]), .A2(a[10]), .B1(n151), .B2(c[10]), .ZN(n13) );
  INV_X1 U24 ( .A(n14), .ZN(carry[12]) );
  AOI22_X1 U25 ( .A1(b[11]), .A2(a[11]), .B1(n152), .B2(c[11]), .ZN(n14) );
  INV_X1 U26 ( .A(n20), .ZN(carry[18]) );
  AOI22_X1 U27 ( .A1(b[17]), .A2(a[17]), .B1(n158), .B2(c[17]), .ZN(n20) );
  INV_X1 U28 ( .A(n25), .ZN(carry[22]) );
  AOI22_X1 U29 ( .A1(b[21]), .A2(a[21]), .B1(n163), .B2(c[21]), .ZN(n25) );
  INV_X1 U30 ( .A(n26), .ZN(carry[23]) );
  AOI22_X1 U31 ( .A1(b[22]), .A2(a[22]), .B1(n164), .B2(c[22]), .ZN(n26) );
  INV_X1 U32 ( .A(n27), .ZN(carry[24]) );
  AOI22_X1 U33 ( .A1(b[23]), .A2(a[23]), .B1(n165), .B2(c[23]), .ZN(n27) );
  INV_X1 U34 ( .A(n29), .ZN(carry[26]) );
  AOI22_X1 U35 ( .A1(b[25]), .A2(a[25]), .B1(n167), .B2(c[25]), .ZN(n29) );
  INV_X1 U36 ( .A(n15), .ZN(carry[13]) );
  AOI22_X1 U37 ( .A1(b[12]), .A2(a[12]), .B1(n153), .B2(c[12]), .ZN(n15) );
  INV_X1 U38 ( .A(n16), .ZN(carry[14]) );
  AOI22_X1 U39 ( .A1(b[13]), .A2(a[13]), .B1(n154), .B2(c[13]), .ZN(n16) );
  INV_X1 U40 ( .A(n17), .ZN(carry[15]) );
  AOI22_X1 U41 ( .A1(b[14]), .A2(a[14]), .B1(n155), .B2(c[14]), .ZN(n17) );
  INV_X1 U42 ( .A(n18), .ZN(carry[16]) );
  AOI22_X1 U43 ( .A1(b[15]), .A2(a[15]), .B1(n156), .B2(c[15]), .ZN(n18) );
  INV_X1 U44 ( .A(n28), .ZN(carry[25]) );
  AOI22_X1 U45 ( .A1(b[24]), .A2(a[24]), .B1(n166), .B2(c[24]), .ZN(n28) );
  INV_X1 U46 ( .A(n31), .ZN(carry[28]) );
  AOI22_X1 U47 ( .A1(b[27]), .A2(a[27]), .B1(n169), .B2(c[27]), .ZN(n31) );
  INV_X1 U48 ( .A(n34), .ZN(carry[30]) );
  AOI22_X1 U49 ( .A1(b[29]), .A2(a[29]), .B1(n171), .B2(c[29]), .ZN(n34) );
  INV_X1 U50 ( .A(n35), .ZN(carry[31]) );
  AOI22_X1 U51 ( .A1(b[30]), .A2(a[30]), .B1(n173), .B2(c[30]), .ZN(n35) );
  INV_X1 U52 ( .A(n36), .ZN(carry[32]) );
  AOI22_X1 U53 ( .A1(b[31]), .A2(a[31]), .B1(n174), .B2(c[31]), .ZN(n36) );
  INV_X1 U54 ( .A(n37), .ZN(carry[33]) );
  AOI22_X1 U55 ( .A1(b[32]), .A2(a[32]), .B1(n175), .B2(c[32]), .ZN(n37) );
  INV_X1 U56 ( .A(n38), .ZN(carry[34]) );
  AOI22_X1 U57 ( .A1(b[33]), .A2(a[33]), .B1(n176), .B2(c[33]), .ZN(n38) );
  INV_X1 U58 ( .A(n147), .ZN(carry[7]) );
  INV_X1 U59 ( .A(n146), .ZN(carry[6]) );
  INV_X1 U60 ( .A(n149), .ZN(carry[9]) );
  INV_X1 U61 ( .A(n12), .ZN(carry[10]) );
  AOI22_X1 U62 ( .A1(b[9]), .A2(a[9]), .B1(n213), .B2(c[9]), .ZN(n12) );
  INV_X1 U63 ( .A(n42), .ZN(carry[38]) );
  AOI22_X1 U64 ( .A1(b[37]), .A2(a[37]), .B1(n180), .B2(c[37]), .ZN(n42) );
  INV_X1 U65 ( .A(n43), .ZN(carry[39]) );
  AOI22_X1 U66 ( .A1(b[38]), .A2(a[38]), .B1(n181), .B2(c[38]), .ZN(n43) );
  INV_X1 U67 ( .A(n45), .ZN(carry[40]) );
  AOI22_X1 U68 ( .A1(b[39]), .A2(a[39]), .B1(n182), .B2(c[39]), .ZN(n45) );
  INV_X1 U69 ( .A(n46), .ZN(carry[41]) );
  AOI22_X1 U70 ( .A1(b[40]), .A2(a[40]), .B1(n184), .B2(c[40]), .ZN(n46) );
  INV_X1 U71 ( .A(n47), .ZN(carry[42]) );
  AOI22_X1 U72 ( .A1(b[41]), .A2(a[41]), .B1(n185), .B2(c[41]), .ZN(n47) );
  INV_X1 U73 ( .A(n40), .ZN(carry[36]) );
  AOI22_X1 U74 ( .A1(b[35]), .A2(a[35]), .B1(n178), .B2(c[35]), .ZN(n40) );
  INV_X1 U75 ( .A(n41), .ZN(carry[37]) );
  AOI22_X1 U76 ( .A1(b[36]), .A2(a[36]), .B1(n179), .B2(c[36]), .ZN(n41) );
  INV_X1 U77 ( .A(n39), .ZN(carry[35]) );
  AOI22_X1 U78 ( .A1(b[34]), .A2(a[34]), .B1(n177), .B2(c[34]), .ZN(n39) );
  INV_X1 U79 ( .A(n60), .ZN(carry[54]) );
  AOI22_X1 U80 ( .A1(b[53]), .A2(a[53]), .B1(n198), .B2(c[53]), .ZN(n60) );
  INV_X1 U81 ( .A(n48), .ZN(carry[43]) );
  AOI22_X1 U82 ( .A1(b[42]), .A2(a[42]), .B1(n186), .B2(c[42]), .ZN(n48) );
  INV_X1 U83 ( .A(n49), .ZN(carry[44]) );
  AOI22_X1 U84 ( .A1(b[43]), .A2(a[43]), .B1(n187), .B2(c[43]), .ZN(n49) );
  INV_X1 U85 ( .A(n50), .ZN(carry[45]) );
  AOI22_X1 U86 ( .A1(b[44]), .A2(a[44]), .B1(n188), .B2(c[44]), .ZN(n50) );
  INV_X1 U87 ( .A(n51), .ZN(carry[46]) );
  AOI22_X1 U88 ( .A1(b[45]), .A2(a[45]), .B1(n189), .B2(c[45]), .ZN(n51) );
  INV_X1 U89 ( .A(n52), .ZN(carry[47]) );
  AOI22_X1 U90 ( .A1(b[46]), .A2(a[46]), .B1(n190), .B2(c[46]), .ZN(n52) );
  INV_X1 U91 ( .A(n53), .ZN(carry[48]) );
  AOI22_X1 U92 ( .A1(b[47]), .A2(a[47]), .B1(n191), .B2(c[47]), .ZN(n53) );
  INV_X1 U93 ( .A(n54), .ZN(carry[49]) );
  AOI22_X1 U94 ( .A1(b[48]), .A2(a[48]), .B1(n192), .B2(c[48]), .ZN(n54) );
  INV_X1 U95 ( .A(n56), .ZN(carry[50]) );
  AOI22_X1 U96 ( .A1(b[49]), .A2(a[49]), .B1(n193), .B2(c[49]), .ZN(n56) );
  INV_X1 U97 ( .A(n57), .ZN(carry[51]) );
  AOI22_X1 U98 ( .A1(b[50]), .A2(a[50]), .B1(n195), .B2(c[50]), .ZN(n57) );
  INV_X1 U99 ( .A(n58), .ZN(carry[52]) );
  AOI22_X1 U100 ( .A1(b[51]), .A2(a[51]), .B1(n196), .B2(c[51]), .ZN(n58) );
  INV_X1 U101 ( .A(n59), .ZN(carry[53]) );
  AOI22_X1 U102 ( .A1(b[52]), .A2(a[52]), .B1(n197), .B2(c[52]), .ZN(n59) );
  INV_X1 U103 ( .A(n61), .ZN(carry[55]) );
  AOI22_X1 U104 ( .A1(b[54]), .A2(a[54]), .B1(n199), .B2(c[54]), .ZN(n61) );
  INV_X1 U105 ( .A(n142), .ZN(carry[60]) );
  AOI22_X1 U106 ( .A1(b[59]), .A2(a[59]), .B1(n204), .B2(c[59]), .ZN(n142) );
  INV_X1 U107 ( .A(n143), .ZN(carry[61]) );
  AOI22_X1 U108 ( .A1(b[60]), .A2(a[60]), .B1(n206), .B2(c[60]), .ZN(n143) );
  INV_X1 U109 ( .A(n144), .ZN(carry[62]) );
  AOI22_X1 U110 ( .A1(b[61]), .A2(a[61]), .B1(n207), .B2(c[61]), .ZN(n144) );
  INV_X1 U111 ( .A(n63), .ZN(carry[57]) );
  AOI22_X1 U112 ( .A1(b[56]), .A2(a[56]), .B1(n201), .B2(c[56]), .ZN(n63) );
  INV_X1 U113 ( .A(n62), .ZN(carry[56]) );
  AOI22_X1 U114 ( .A1(b[55]), .A2(a[55]), .B1(n200), .B2(c[55]), .ZN(n62) );
  INV_X1 U115 ( .A(n139), .ZN(carry[58]) );
  AOI22_X1 U116 ( .A1(b[57]), .A2(a[57]), .B1(n202), .B2(c[57]), .ZN(n139) );
  INV_X1 U117 ( .A(n140), .ZN(carry[59]) );
  AOI22_X1 U118 ( .A1(b[58]), .A2(a[58]), .B1(n203), .B2(c[58]), .ZN(n140) );
  INV_X1 U119 ( .A(n145), .ZN(carry[63]) );
  AOI22_X1 U120 ( .A1(b[62]), .A2(a[62]), .B1(n208), .B2(c[62]), .ZN(n145) );
  INV_X1 U121 ( .A(n148), .ZN(carry[8]) );
  INV_X1 U122 ( .A(n141), .ZN(carry[5]) );
  INV_X1 U123 ( .A(n22), .ZN(carry[1]) );
  AOI22_X1 U124 ( .A1(b[0]), .A2(a[0]), .B1(n150), .B2(c[0]), .ZN(n22) );
  INV_X1 U125 ( .A(n33), .ZN(carry[2]) );
  AOI22_X1 U126 ( .A1(b[1]), .A2(a[1]), .B1(n161), .B2(c[1]), .ZN(n33) );
  INV_X1 U127 ( .A(n44), .ZN(carry[3]) );
  AOI22_X1 U129 ( .A1(b[2]), .A2(a[2]), .B1(n172), .B2(c[2]), .ZN(n44) );
  INV_X1 U148 ( .A(n55), .ZN(carry[4]) );
  AOI22_X1 U254 ( .A1(b[3]), .A2(a[3]), .B1(n183), .B2(c[3]), .ZN(n55) );
  NAND2_X1 U256 ( .A1(c[8]), .A2(n8), .ZN(n9) );
  NAND2_X1 U257 ( .A1(n212), .A2(n7), .ZN(n10) );
  NAND2_X1 U258 ( .A1(n9), .A2(n10), .ZN(result[8]) );
  INV_X1 U259 ( .A(c[8]), .ZN(n7) );
  INV_X1 U260 ( .A(n212), .ZN(n8) );
  CLKBUF_X1 U261 ( .A(b[5]), .Z(n11) );
  AOI22_X1 U262 ( .A1(b[4]), .A2(a[4]), .B1(n194), .B2(c[4]), .ZN(n141) );
  AOI22_X1 U263 ( .A1(b[6]), .A2(a[6]), .B1(n210), .B2(c[6]), .ZN(n147) );
  AOI22_X1 U264 ( .A1(b[8]), .A2(a[8]), .B1(n212), .B2(c[8]), .ZN(n149) );
  AOI22_X1 U265 ( .A1(n11), .A2(n5), .B1(n205), .B2(c[5]), .ZN(n146) );
  AOI22_X1 U266 ( .A1(b[7]), .A2(a[7]), .B1(c[7]), .B2(n211), .ZN(n148) );
endmodule


module TM ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;
  wire   shiftedA_7__63_, shiftedA_7__37_, shiftedA_7__36_, shiftedA_7__35_,
         shiftedA_7__34_, shiftedA_7__33_, shiftedA_7__32_, shiftedA_7__31_,
         shiftedA_7__30_, shiftedA_7__29_, shiftedA_7__28_, shiftedA_7__27_,
         shiftedA_7__26_, shiftedA_7__25_, shiftedA_7__24_, shiftedA_7__23_,
         shiftedA_7__22_, shiftedA_7__21_, shiftedA_7__20_, shiftedA_7__19_,
         shiftedA_7__18_, shiftedA_7__17_, shiftedA_7__16_, shiftedA_7__15_,
         shiftedA_7__14_, shiftedA_7__13_, shiftedA_7__12_, shiftedA_7__11_,
         shiftedA_7__10_, shiftedA_7__9_, shiftedA_7__8_, shiftedA_7__7_,
         shiftedA_6__63_, shiftedA_6__36_, shiftedA_6__35_, shiftedA_6__34_,
         shiftedA_6__33_, shiftedA_6__32_, shiftedA_6__31_, shiftedA_6__30_,
         shiftedA_6__29_, shiftedA_6__28_, shiftedA_6__27_, shiftedA_6__26_,
         shiftedA_6__25_, shiftedA_6__24_, shiftedA_6__23_, shiftedA_6__22_,
         shiftedA_6__21_, shiftedA_6__20_, shiftedA_6__19_, shiftedA_6__18_,
         shiftedA_6__17_, shiftedA_6__16_, shiftedA_6__15_, shiftedA_6__14_,
         shiftedA_6__13_, shiftedA_6__12_, shiftedA_6__11_, shiftedA_6__10_,
         shiftedA_6__9_, shiftedA_6__8_, shiftedA_6__7_, shiftedA_6__6_,
         shiftedA_5__63_, shiftedA_5__35_, shiftedA_5__34_, shiftedA_5__33_,
         shiftedA_5__32_, shiftedA_5__31_, shiftedA_5__30_, shiftedA_5__29_,
         shiftedA_5__28_, shiftedA_5__27_, shiftedA_5__26_, shiftedA_5__25_,
         shiftedA_5__24_, shiftedA_5__23_, shiftedA_5__22_, shiftedA_5__21_,
         shiftedA_5__20_, shiftedA_5__19_, shiftedA_5__18_, shiftedA_5__17_,
         shiftedA_5__16_, shiftedA_5__15_, shiftedA_5__14_, shiftedA_5__13_,
         shiftedA_5__12_, shiftedA_5__11_, shiftedA_5__10_, shiftedA_5__9_,
         shiftedA_5__8_, shiftedA_5__7_, shiftedA_5__6_, shiftedA_5__5_,
         shiftedA_4__63_, shiftedA_4__34_, shiftedA_4__33_, shiftedA_4__32_,
         shiftedA_4__31_, shiftedA_4__30_, shiftedA_4__29_, shiftedA_4__28_,
         shiftedA_4__27_, shiftedA_4__26_, shiftedA_4__25_, shiftedA_4__24_,
         shiftedA_4__23_, shiftedA_4__22_, shiftedA_4__21_, shiftedA_4__20_,
         shiftedA_4__19_, shiftedA_4__18_, shiftedA_4__17_, shiftedA_4__16_,
         shiftedA_4__15_, shiftedA_4__14_, shiftedA_4__13_, shiftedA_4__12_,
         shiftedA_4__11_, shiftedA_4__10_, shiftedA_4__9_, shiftedA_4__8_,
         shiftedA_4__7_, shiftedA_4__6_, shiftedA_4__5_, shiftedA_4__4_,
         shiftedA_3__63_, shiftedA_3__33_, shiftedA_3__32_, shiftedA_3__31_,
         shiftedA_3__30_, shiftedA_3__29_, shiftedA_3__28_, shiftedA_3__27_,
         shiftedA_3__26_, shiftedA_3__25_, shiftedA_3__24_, shiftedA_3__23_,
         shiftedA_3__22_, shiftedA_3__21_, shiftedA_3__20_, shiftedA_3__19_,
         shiftedA_3__18_, shiftedA_3__17_, shiftedA_3__16_, shiftedA_3__15_,
         shiftedA_3__14_, shiftedA_3__13_, shiftedA_3__12_, shiftedA_3__11_,
         shiftedA_3__10_, shiftedA_3__9_, shiftedA_3__8_, shiftedA_3__7_,
         shiftedA_3__6_, shiftedA_3__5_, shiftedA_3__4_, shiftedA_3__3_,
         shiftedA_2__63_, shiftedA_2__32_, shiftedA_2__31_, shiftedA_2__30_,
         shiftedA_2__29_, shiftedA_2__28_, shiftedA_2__27_, shiftedA_2__26_,
         shiftedA_2__25_, shiftedA_2__24_, shiftedA_2__23_, shiftedA_2__22_,
         shiftedA_2__21_, shiftedA_2__20_, shiftedA_2__19_, shiftedA_2__18_,
         shiftedA_2__17_, shiftedA_2__16_, shiftedA_2__15_, shiftedA_2__14_,
         shiftedA_2__13_, shiftedA_2__12_, shiftedA_2__11_, shiftedA_2__10_,
         shiftedA_2__9_, shiftedA_2__8_, shiftedA_2__7_, shiftedA_2__6_,
         shiftedA_2__5_, shiftedA_2__4_, shiftedA_2__3_, shiftedA_2__2_,
         shiftedA_1__63_, shiftedA_1__31_, shiftedA_1__30_, shiftedA_1__29_,
         shiftedA_1__28_, shiftedA_1__27_, shiftedA_1__26_, shiftedA_1__25_,
         shiftedA_1__24_, shiftedA_1__23_, shiftedA_1__22_, shiftedA_1__21_,
         shiftedA_1__20_, shiftedA_1__19_, shiftedA_1__18_, shiftedA_1__17_,
         shiftedA_1__16_, shiftedA_1__15_, shiftedA_1__14_, shiftedA_1__13_,
         shiftedA_1__12_, shiftedA_1__11_, shiftedA_1__10_, shiftedA_1__9_,
         shiftedA_1__8_, shiftedA_1__7_, shiftedA_1__6_, shiftedA_1__5_,
         shiftedA_1__4_, shiftedA_1__3_, shiftedA_1__2_, shiftedA_1__1_,
         shiftedA_0__63_, shiftedA_0__30_, shiftedA_0__29_, shiftedA_0__28_,
         shiftedA_0__27_, shiftedA_0__26_, shiftedA_0__25_, shiftedA_0__24_,
         shiftedA_0__23_, shiftedA_0__22_, shiftedA_0__21_, shiftedA_0__20_,
         shiftedA_0__19_, shiftedA_0__18_, shiftedA_0__17_, shiftedA_0__16_,
         shiftedA_0__15_, shiftedA_0__14_, shiftedA_0__13_, shiftedA_0__12_,
         shiftedA_0__11_, shiftedA_0__10_, shiftedA_0__9_, shiftedA_0__8_,
         shiftedA_0__7_, shiftedA_0__6_, shiftedA_0__5_, shiftedA_0__4_,
         shiftedA_0__3_, shiftedA_0__2_, shiftedA_0__1_, shiftedA_0__0_,
         shiftedA_63__63_, shiftedA_62__63_, shiftedA_61__63_,
         shiftedA_60__63_, shiftedA_59__63_, shiftedA_58__63_,
         shiftedA_57__63_, shiftedA_56__63_, shiftedA_55__63_,
         shiftedA_54__63_, shiftedA_53__63_, shiftedA_52__63_,
         shiftedA_51__63_, shiftedA_50__63_, shiftedA_49__63_,
         shiftedA_48__63_, shiftedA_47__63_, shiftedA_46__63_,
         shiftedA_45__63_, shiftedA_44__63_, shiftedA_43__63_,
         shiftedA_42__63_, shiftedA_41__63_, shiftedA_40__63_,
         shiftedA_39__63_, shiftedA_38__63_, shiftedA_37__63_,
         shiftedA_36__63_, shiftedA_35__63_, shiftedA_34__63_,
         shiftedA_33__63_, shiftedA_32__63_, shiftedA_30__63_,
         shiftedA_30__60_, shiftedA_30__59_, shiftedA_30__58_,
         shiftedA_30__57_, shiftedA_30__56_, shiftedA_30__55_,
         shiftedA_30__54_, shiftedA_30__53_, shiftedA_30__52_,
         shiftedA_30__51_, shiftedA_30__50_, shiftedA_30__49_,
         shiftedA_30__48_, shiftedA_30__47_, shiftedA_30__46_,
         shiftedA_30__45_, shiftedA_30__44_, shiftedA_30__43_,
         shiftedA_30__42_, shiftedA_30__41_, shiftedA_30__40_,
         shiftedA_30__39_, shiftedA_30__38_, shiftedA_30__37_,
         shiftedA_30__36_, shiftedA_30__35_, shiftedA_30__34_,
         shiftedA_30__33_, shiftedA_30__32_, shiftedA_30__31_,
         shiftedA_30__30_, shiftedA_29__63_, shiftedA_29__59_,
         shiftedA_29__58_, shiftedA_29__57_, shiftedA_29__56_,
         shiftedA_29__55_, shiftedA_29__54_, shiftedA_29__53_,
         shiftedA_29__52_, shiftedA_29__51_, shiftedA_29__50_,
         shiftedA_29__49_, shiftedA_29__48_, shiftedA_29__47_,
         shiftedA_29__46_, shiftedA_29__45_, shiftedA_29__44_,
         shiftedA_29__43_, shiftedA_29__42_, shiftedA_29__41_,
         shiftedA_29__40_, shiftedA_29__39_, shiftedA_29__38_,
         shiftedA_29__37_, shiftedA_29__36_, shiftedA_29__35_,
         shiftedA_29__34_, shiftedA_29__33_, shiftedA_29__32_,
         shiftedA_29__31_, shiftedA_29__30_, shiftedA_29__29_,
         shiftedA_28__63_, shiftedA_28__58_, shiftedA_28__57_,
         shiftedA_28__56_, shiftedA_28__55_, shiftedA_28__54_,
         shiftedA_28__53_, shiftedA_28__52_, shiftedA_28__51_,
         shiftedA_28__50_, shiftedA_28__49_, shiftedA_28__48_,
         shiftedA_28__47_, shiftedA_28__46_, shiftedA_28__45_,
         shiftedA_28__44_, shiftedA_28__43_, shiftedA_28__42_,
         shiftedA_28__41_, shiftedA_28__40_, shiftedA_28__39_,
         shiftedA_28__38_, shiftedA_28__37_, shiftedA_28__36_,
         shiftedA_28__35_, shiftedA_28__34_, shiftedA_28__33_,
         shiftedA_28__32_, shiftedA_28__31_, shiftedA_28__30_,
         shiftedA_28__29_, shiftedA_28__28_, shiftedA_27__63_,
         shiftedA_27__57_, shiftedA_27__56_, shiftedA_27__55_,
         shiftedA_27__54_, shiftedA_27__53_, shiftedA_27__52_,
         shiftedA_27__51_, shiftedA_27__50_, shiftedA_27__49_,
         shiftedA_27__48_, shiftedA_27__47_, shiftedA_27__46_,
         shiftedA_27__45_, shiftedA_27__44_, shiftedA_27__43_,
         shiftedA_27__42_, shiftedA_27__41_, shiftedA_27__40_,
         shiftedA_27__39_, shiftedA_27__38_, shiftedA_27__37_,
         shiftedA_27__36_, shiftedA_27__35_, shiftedA_27__34_,
         shiftedA_27__33_, shiftedA_27__32_, shiftedA_27__31_,
         shiftedA_27__30_, shiftedA_27__29_, shiftedA_27__28_,
         shiftedA_27__27_, shiftedA_26__63_, shiftedA_26__56_,
         shiftedA_26__55_, shiftedA_26__54_, shiftedA_26__53_,
         shiftedA_26__52_, shiftedA_26__51_, shiftedA_26__50_,
         shiftedA_26__49_, shiftedA_26__48_, shiftedA_26__47_,
         shiftedA_26__46_, shiftedA_26__45_, shiftedA_26__44_,
         shiftedA_26__43_, shiftedA_26__42_, shiftedA_26__41_,
         shiftedA_26__40_, shiftedA_26__39_, shiftedA_26__38_,
         shiftedA_26__37_, shiftedA_26__36_, shiftedA_26__35_,
         shiftedA_26__34_, shiftedA_26__33_, shiftedA_26__32_,
         shiftedA_26__31_, shiftedA_26__30_, shiftedA_26__29_,
         shiftedA_26__28_, shiftedA_26__27_, shiftedA_26__26_,
         shiftedA_25__63_, shiftedA_25__55_, shiftedA_25__54_,
         shiftedA_25__53_, shiftedA_25__52_, shiftedA_25__51_,
         shiftedA_25__50_, shiftedA_25__49_, shiftedA_25__48_,
         shiftedA_25__47_, shiftedA_25__46_, shiftedA_25__45_,
         shiftedA_25__44_, shiftedA_25__43_, shiftedA_25__42_,
         shiftedA_25__41_, shiftedA_25__40_, shiftedA_25__39_,
         shiftedA_25__38_, shiftedA_25__37_, shiftedA_25__36_,
         shiftedA_25__35_, shiftedA_25__34_, shiftedA_25__33_,
         shiftedA_25__32_, shiftedA_25__31_, shiftedA_25__30_,
         shiftedA_25__29_, shiftedA_25__28_, shiftedA_25__27_,
         shiftedA_25__26_, shiftedA_25__25_, shiftedA_24__63_,
         shiftedA_24__54_, shiftedA_24__53_, shiftedA_24__52_,
         shiftedA_24__51_, shiftedA_24__50_, shiftedA_24__49_,
         shiftedA_24__48_, shiftedA_24__47_, shiftedA_24__46_,
         shiftedA_24__45_, shiftedA_24__44_, shiftedA_24__43_,
         shiftedA_24__42_, shiftedA_24__41_, shiftedA_24__40_,
         shiftedA_24__39_, shiftedA_24__38_, shiftedA_24__37_,
         shiftedA_24__36_, shiftedA_24__35_, shiftedA_24__34_,
         shiftedA_24__33_, shiftedA_24__32_, shiftedA_24__31_,
         shiftedA_24__30_, shiftedA_24__29_, shiftedA_24__28_,
         shiftedA_24__27_, shiftedA_24__26_, shiftedA_24__25_,
         shiftedA_24__24_, shiftedA_23__63_, shiftedA_23__53_,
         shiftedA_23__52_, shiftedA_23__51_, shiftedA_23__50_,
         shiftedA_23__49_, shiftedA_23__48_, shiftedA_23__47_,
         shiftedA_23__46_, shiftedA_23__45_, shiftedA_23__44_,
         shiftedA_23__43_, shiftedA_23__42_, shiftedA_23__41_,
         shiftedA_23__40_, shiftedA_23__39_, shiftedA_23__38_,
         shiftedA_23__37_, shiftedA_23__36_, shiftedA_23__35_,
         shiftedA_23__34_, shiftedA_23__33_, shiftedA_23__32_,
         shiftedA_23__31_, shiftedA_23__30_, shiftedA_23__29_,
         shiftedA_23__28_, shiftedA_23__27_, shiftedA_23__26_,
         shiftedA_23__25_, shiftedA_23__24_, shiftedA_23__23_,
         shiftedA_22__63_, shiftedA_22__52_, shiftedA_22__51_,
         shiftedA_22__50_, shiftedA_22__49_, shiftedA_22__48_,
         shiftedA_22__47_, shiftedA_22__46_, shiftedA_22__45_,
         shiftedA_22__44_, shiftedA_22__43_, shiftedA_22__42_,
         shiftedA_22__41_, shiftedA_22__40_, shiftedA_22__39_,
         shiftedA_22__38_, shiftedA_22__37_, shiftedA_22__36_,
         shiftedA_22__35_, shiftedA_22__34_, shiftedA_22__33_,
         shiftedA_22__32_, shiftedA_22__31_, shiftedA_22__30_,
         shiftedA_22__29_, shiftedA_22__28_, shiftedA_22__27_,
         shiftedA_22__26_, shiftedA_22__25_, shiftedA_22__24_,
         shiftedA_22__23_, shiftedA_22__22_, shiftedA_21__63_,
         shiftedA_21__51_, shiftedA_21__50_, shiftedA_21__49_,
         shiftedA_21__48_, shiftedA_21__47_, shiftedA_21__46_,
         shiftedA_21__45_, shiftedA_21__44_, shiftedA_21__43_,
         shiftedA_21__42_, shiftedA_21__41_, shiftedA_21__40_,
         shiftedA_21__39_, shiftedA_21__38_, shiftedA_21__37_,
         shiftedA_21__36_, shiftedA_21__35_, shiftedA_21__34_,
         shiftedA_21__33_, shiftedA_21__32_, shiftedA_21__31_,
         shiftedA_21__30_, shiftedA_21__29_, shiftedA_21__28_,
         shiftedA_21__27_, shiftedA_21__26_, shiftedA_21__25_,
         shiftedA_21__24_, shiftedA_21__23_, shiftedA_21__22_,
         shiftedA_21__21_, shiftedA_20__63_, shiftedA_20__50_,
         shiftedA_20__49_, shiftedA_20__48_, shiftedA_20__47_,
         shiftedA_20__46_, shiftedA_20__45_, shiftedA_20__44_,
         shiftedA_20__43_, shiftedA_20__42_, shiftedA_20__41_,
         shiftedA_20__40_, shiftedA_20__39_, shiftedA_20__38_,
         shiftedA_20__37_, shiftedA_20__36_, shiftedA_20__35_,
         shiftedA_20__34_, shiftedA_20__33_, shiftedA_20__32_,
         shiftedA_20__31_, shiftedA_20__30_, shiftedA_20__29_,
         shiftedA_20__28_, shiftedA_20__27_, shiftedA_20__26_,
         shiftedA_20__25_, shiftedA_20__24_, shiftedA_20__23_,
         shiftedA_20__22_, shiftedA_20__21_, shiftedA_20__20_,
         shiftedA_19__63_, shiftedA_19__49_, shiftedA_19__48_,
         shiftedA_19__47_, shiftedA_19__46_, shiftedA_19__45_,
         shiftedA_19__44_, shiftedA_19__43_, shiftedA_19__42_,
         shiftedA_19__41_, shiftedA_19__40_, shiftedA_19__39_,
         shiftedA_19__38_, shiftedA_19__37_, shiftedA_19__36_,
         shiftedA_19__35_, shiftedA_19__34_, shiftedA_19__33_,
         shiftedA_19__32_, shiftedA_19__31_, shiftedA_19__30_,
         shiftedA_19__29_, shiftedA_19__28_, shiftedA_19__27_,
         shiftedA_19__26_, shiftedA_19__25_, shiftedA_19__24_,
         shiftedA_19__23_, shiftedA_19__22_, shiftedA_19__21_,
         shiftedA_19__20_, shiftedA_19__19_, shiftedA_18__63_,
         shiftedA_18__48_, shiftedA_18__47_, shiftedA_18__46_,
         shiftedA_18__45_, shiftedA_18__44_, shiftedA_18__43_,
         shiftedA_18__42_, shiftedA_18__41_, shiftedA_18__40_,
         shiftedA_18__39_, shiftedA_18__38_, shiftedA_18__37_,
         shiftedA_18__36_, shiftedA_18__35_, shiftedA_18__34_,
         shiftedA_18__33_, shiftedA_18__32_, shiftedA_18__31_,
         shiftedA_18__30_, shiftedA_18__29_, shiftedA_18__28_,
         shiftedA_18__27_, shiftedA_18__26_, shiftedA_18__25_,
         shiftedA_18__24_, shiftedA_18__23_, shiftedA_18__22_,
         shiftedA_18__21_, shiftedA_18__20_, shiftedA_18__19_,
         shiftedA_18__18_, shiftedA_17__63_, shiftedA_17__47_,
         shiftedA_17__46_, shiftedA_17__45_, shiftedA_17__44_,
         shiftedA_17__43_, shiftedA_17__42_, shiftedA_17__41_,
         shiftedA_17__40_, shiftedA_17__39_, shiftedA_17__38_,
         shiftedA_17__37_, shiftedA_17__36_, shiftedA_17__35_,
         shiftedA_17__34_, shiftedA_17__33_, shiftedA_17__32_,
         shiftedA_17__31_, shiftedA_17__30_, shiftedA_17__29_,
         shiftedA_17__28_, shiftedA_17__27_, shiftedA_17__26_,
         shiftedA_17__25_, shiftedA_17__24_, shiftedA_17__23_,
         shiftedA_17__22_, shiftedA_17__21_, shiftedA_17__20_,
         shiftedA_17__19_, shiftedA_17__18_, shiftedA_17__17_,
         shiftedA_16__63_, shiftedA_16__46_, shiftedA_16__45_,
         shiftedA_16__44_, shiftedA_16__43_, shiftedA_16__42_,
         shiftedA_16__41_, shiftedA_16__40_, shiftedA_16__39_,
         shiftedA_16__38_, shiftedA_16__37_, shiftedA_16__36_,
         shiftedA_16__35_, shiftedA_16__34_, shiftedA_16__33_,
         shiftedA_16__32_, shiftedA_16__31_, shiftedA_16__30_,
         shiftedA_16__29_, shiftedA_16__28_, shiftedA_16__27_,
         shiftedA_16__26_, shiftedA_16__25_, shiftedA_16__24_,
         shiftedA_16__23_, shiftedA_16__22_, shiftedA_16__21_,
         shiftedA_16__20_, shiftedA_16__19_, shiftedA_16__18_,
         shiftedA_16__17_, shiftedA_16__16_, shiftedA_15__63_,
         shiftedA_15__45_, shiftedA_15__44_, shiftedA_15__43_,
         shiftedA_15__42_, shiftedA_15__41_, shiftedA_15__40_,
         shiftedA_15__39_, shiftedA_15__38_, shiftedA_15__37_,
         shiftedA_15__36_, shiftedA_15__35_, shiftedA_15__34_,
         shiftedA_15__33_, shiftedA_15__32_, shiftedA_15__31_,
         shiftedA_15__30_, shiftedA_15__29_, shiftedA_15__28_,
         shiftedA_15__27_, shiftedA_15__26_, shiftedA_15__25_,
         shiftedA_15__24_, shiftedA_15__23_, shiftedA_15__22_,
         shiftedA_15__21_, shiftedA_15__20_, shiftedA_15__19_,
         shiftedA_15__18_, shiftedA_15__17_, shiftedA_15__16_,
         shiftedA_15__15_, shiftedA_14__63_, shiftedA_14__44_,
         shiftedA_14__43_, shiftedA_14__42_, shiftedA_14__41_,
         shiftedA_14__40_, shiftedA_14__39_, shiftedA_14__38_,
         shiftedA_14__37_, shiftedA_14__36_, shiftedA_14__35_,
         shiftedA_14__34_, shiftedA_14__33_, shiftedA_14__32_,
         shiftedA_14__31_, shiftedA_14__30_, shiftedA_14__29_,
         shiftedA_14__28_, shiftedA_14__27_, shiftedA_14__26_,
         shiftedA_14__25_, shiftedA_14__24_, shiftedA_14__23_,
         shiftedA_14__22_, shiftedA_14__21_, shiftedA_14__20_,
         shiftedA_14__19_, shiftedA_14__18_, shiftedA_14__17_,
         shiftedA_14__16_, shiftedA_14__15_, shiftedA_14__14_,
         shiftedA_13__63_, shiftedA_13__43_, shiftedA_13__42_,
         shiftedA_13__41_, shiftedA_13__40_, shiftedA_13__39_,
         shiftedA_13__38_, shiftedA_13__37_, shiftedA_13__36_,
         shiftedA_13__35_, shiftedA_13__34_, shiftedA_13__33_,
         shiftedA_13__32_, shiftedA_13__31_, shiftedA_13__30_,
         shiftedA_13__29_, shiftedA_13__28_, shiftedA_13__27_,
         shiftedA_13__26_, shiftedA_13__25_, shiftedA_13__24_,
         shiftedA_13__23_, shiftedA_13__22_, shiftedA_13__21_,
         shiftedA_13__20_, shiftedA_13__19_, shiftedA_13__18_,
         shiftedA_13__17_, shiftedA_13__16_, shiftedA_13__15_,
         shiftedA_13__14_, shiftedA_13__13_, shiftedA_12__63_,
         shiftedA_12__42_, shiftedA_12__41_, shiftedA_12__40_,
         shiftedA_12__39_, shiftedA_12__38_, shiftedA_12__37_,
         shiftedA_12__36_, shiftedA_12__35_, shiftedA_12__34_,
         shiftedA_12__33_, shiftedA_12__32_, shiftedA_12__31_,
         shiftedA_12__30_, shiftedA_12__29_, shiftedA_12__28_,
         shiftedA_12__27_, shiftedA_12__26_, shiftedA_12__25_,
         shiftedA_12__24_, shiftedA_12__23_, shiftedA_12__22_,
         shiftedA_12__21_, shiftedA_12__20_, shiftedA_12__19_,
         shiftedA_12__18_, shiftedA_12__17_, shiftedA_12__16_,
         shiftedA_12__15_, shiftedA_12__14_, shiftedA_12__13_,
         shiftedA_12__12_, shiftedA_11__63_, shiftedA_11__41_,
         shiftedA_11__40_, shiftedA_11__39_, shiftedA_11__38_,
         shiftedA_11__37_, shiftedA_11__36_, shiftedA_11__35_,
         shiftedA_11__34_, shiftedA_11__33_, shiftedA_11__32_,
         shiftedA_11__31_, shiftedA_11__30_, shiftedA_11__29_,
         shiftedA_11__28_, shiftedA_11__27_, shiftedA_11__26_,
         shiftedA_11__25_, shiftedA_11__24_, shiftedA_11__23_,
         shiftedA_11__22_, shiftedA_11__21_, shiftedA_11__20_,
         shiftedA_11__19_, shiftedA_11__18_, shiftedA_11__17_,
         shiftedA_11__16_, shiftedA_11__15_, shiftedA_11__14_,
         shiftedA_11__13_, shiftedA_11__12_, shiftedA_11__11_,
         shiftedA_10__63_, shiftedA_10__40_, shiftedA_10__39_,
         shiftedA_10__38_, shiftedA_10__37_, shiftedA_10__36_,
         shiftedA_10__35_, shiftedA_10__34_, shiftedA_10__33_,
         shiftedA_10__32_, shiftedA_10__31_, shiftedA_10__30_,
         shiftedA_10__29_, shiftedA_10__28_, shiftedA_10__27_,
         shiftedA_10__26_, shiftedA_10__25_, shiftedA_10__24_,
         shiftedA_10__23_, shiftedA_10__22_, shiftedA_10__21_,
         shiftedA_10__20_, shiftedA_10__19_, shiftedA_10__18_,
         shiftedA_10__17_, shiftedA_10__16_, shiftedA_10__15_,
         shiftedA_10__14_, shiftedA_10__13_, shiftedA_10__12_,
         shiftedA_10__11_, shiftedA_10__10_, shiftedA_9__63_, shiftedA_9__39_,
         shiftedA_9__38_, shiftedA_9__37_, shiftedA_9__36_, shiftedA_9__35_,
         shiftedA_9__34_, shiftedA_9__33_, shiftedA_9__32_, shiftedA_9__31_,
         shiftedA_9__30_, shiftedA_9__29_, shiftedA_9__28_, shiftedA_9__27_,
         shiftedA_9__26_, shiftedA_9__25_, shiftedA_9__24_, shiftedA_9__23_,
         shiftedA_9__22_, shiftedA_9__21_, shiftedA_9__20_, shiftedA_9__19_,
         shiftedA_9__18_, shiftedA_9__17_, shiftedA_9__16_, shiftedA_9__15_,
         shiftedA_9__14_, shiftedA_9__13_, shiftedA_9__12_, shiftedA_9__11_,
         shiftedA_9__10_, shiftedA_9__9_, shiftedA_8__63_, shiftedA_8__38_,
         shiftedA_8__37_, shiftedA_8__36_, shiftedA_8__35_, shiftedA_8__34_,
         shiftedA_8__33_, shiftedA_8__32_, shiftedA_8__31_, shiftedA_8__30_,
         shiftedA_8__29_, shiftedA_8__28_, shiftedA_8__27_, shiftedA_8__26_,
         shiftedA_8__25_, shiftedA_8__24_, shiftedA_8__23_, shiftedA_8__22_,
         shiftedA_8__21_, shiftedA_8__20_, shiftedA_8__19_, shiftedA_8__18_,
         shiftedA_8__17_, shiftedA_8__16_, shiftedA_8__15_, shiftedA_8__14_,
         shiftedA_8__13_, shiftedA_8__12_, shiftedA_8__11_, shiftedA_8__10_,
         shiftedA_8__9_, shiftedA_8__8_, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n27, n28, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n26, n29, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375;
  wire   [1343:0] adderResult_level1;
  wire   [1343:0] carry_level1;
  wire   [895:0] adderResult_level2;
  wire   [895:0] carry_level2;
  wire   [575:0] adderResult_level3;
  wire   [575:0] carry_level3;
  wire   [383:0] adderResult_level4;
  wire   [383:0] carry_level4;
  wire   [255:0] adderResult_level5;
  wire   [255:0] carry_level5;
  wire   [191:0] adderResult_level6;
  wire   [191:0] carry_level6;
  wire   [127:0] adderResult_level7;
  wire   [127:0] carry_level7;
  wire   [63:0] adderResult_level8;
  wire   [63:0] carry_level8;
  wire   [63:0] adderResult_level9;
  wire   [63:0] carry_level9;
  wire   [63:0] adderResult_level10;
  wire   [63:0] carry_level10;

  BWAdder_0 level1_0__adder ( .a({n348, n348, n348, n348, n348, n348, n348, 
        n348, n348, n347, n347, n347, n347, n347, n347, n347, n347, n347, n347, 
        n347, n347, n346, n346, n346, n346, n346, n346, n346, n346, n346, n346, 
        n346, n346, shiftedA_0__30_, shiftedA_0__29_, shiftedA_0__28_, 
        shiftedA_0__27_, shiftedA_0__26_, shiftedA_0__25_, shiftedA_0__24_, 
        shiftedA_0__23_, shiftedA_0__22_, shiftedA_0__21_, shiftedA_0__20_, 
        shiftedA_0__19_, shiftedA_0__18_, shiftedA_0__17_, shiftedA_0__16_, 
        shiftedA_0__15_, shiftedA_0__14_, shiftedA_0__13_, shiftedA_0__12_, 
        shiftedA_0__11_, shiftedA_0__10_, shiftedA_0__9_, shiftedA_0__8_, 
        shiftedA_0__7_, shiftedA_0__6_, shiftedA_0__5_, shiftedA_0__4_, 
        shiftedA_0__3_, shiftedA_0__2_, shiftedA_0__1_, shiftedA_0__0_}), .b({
        n351, n351, n351, n351, n351, n351, n351, n351, n350, n350, n350, n350, 
        n350, n350, n350, n350, n350, n350, n350, n350, n349, n349, n349, n349, 
        n349, n349, n349, n349, n349, n349, n349, n349, shiftedA_1__31_, 
        shiftedA_1__30_, shiftedA_1__29_, shiftedA_1__28_, shiftedA_1__27_, 
        shiftedA_1__26_, shiftedA_1__25_, shiftedA_1__24_, shiftedA_1__23_, 
        shiftedA_1__22_, shiftedA_1__21_, shiftedA_1__20_, shiftedA_1__19_, 
        shiftedA_1__18_, shiftedA_1__17_, shiftedA_1__16_, shiftedA_1__15_, 
        shiftedA_1__14_, shiftedA_1__13_, shiftedA_1__12_, shiftedA_1__11_, 
        shiftedA_1__10_, shiftedA_1__9_, shiftedA_1__8_, shiftedA_1__7_, 
        shiftedA_1__6_, shiftedA_1__5_, shiftedA_1__4_, shiftedA_1__3_, 
        shiftedA_1__2_, shiftedA_1__1_, 1'b0}), .c({n354, n354, n354, n354, 
        n354, n354, n354, n353, n353, n353, n353, n353, n353, n353, n353, n353, 
        n353, n353, n353, n352, n352, n352, n352, n352, n352, n352, n352, n352, 
        n352, n352, n352, shiftedA_2__32_, shiftedA_2__31_, shiftedA_2__30_, 
        shiftedA_2__29_, shiftedA_2__28_, shiftedA_2__27_, shiftedA_2__26_, 
        shiftedA_2__25_, shiftedA_2__24_, shiftedA_2__23_, shiftedA_2__22_, 
        shiftedA_2__21_, shiftedA_2__20_, shiftedA_2__19_, shiftedA_2__18_, 
        shiftedA_2__17_, shiftedA_2__16_, shiftedA_2__15_, shiftedA_2__14_, 
        shiftedA_2__13_, shiftedA_2__12_, shiftedA_2__11_, shiftedA_2__10_, 
        shiftedA_2__9_, shiftedA_2__8_, shiftedA_2__7_, shiftedA_2__6_, 
        shiftedA_2__5_, shiftedA_2__4_, shiftedA_2__3_, shiftedA_2__2_, 1'b0, 
        1'b0}), .result(adderResult_level1[63:0]), .carry(carry_level1[63:0])
         );
  BWAdder_61 level1_1__adder ( .a({n357, n357, n357, n357, n357, n357, n356, 
        n356, n356, n356, n356, n356, n356, n356, n356, n356, n356, n356, n355, 
        n355, n355, n355, n355, n355, n355, n355, n355, n355, n355, n355, 
        shiftedA_3__33_, shiftedA_3__32_, shiftedA_3__31_, shiftedA_3__30_, 
        shiftedA_3__29_, shiftedA_3__28_, shiftedA_3__27_, shiftedA_3__26_, 
        shiftedA_3__25_, shiftedA_3__24_, shiftedA_3__23_, shiftedA_3__22_, 
        shiftedA_3__21_, shiftedA_3__20_, shiftedA_3__19_, shiftedA_3__18_, 
        shiftedA_3__17_, shiftedA_3__16_, shiftedA_3__15_, shiftedA_3__14_, 
        shiftedA_3__13_, shiftedA_3__12_, shiftedA_3__11_, shiftedA_3__10_, 
        shiftedA_3__9_, shiftedA_3__8_, shiftedA_3__7_, shiftedA_3__6_, 
        shiftedA_3__5_, shiftedA_3__4_, shiftedA_3__3_, 1'b0, 1'b0, 1'b0}), 
        .b({n360, n360, n360, n360, n360, n359, n359, n359, n359, n359, n359, 
        n359, n359, n359, n359, n359, n359, n358, n358, n358, n358, n358, n358, 
        n358, n358, n358, n358, n358, n358, shiftedA_4__34_, shiftedA_4__33_, 
        shiftedA_4__32_, shiftedA_4__31_, shiftedA_4__30_, shiftedA_4__29_, 
        shiftedA_4__28_, shiftedA_4__27_, shiftedA_4__26_, shiftedA_4__25_, 
        shiftedA_4__24_, shiftedA_4__23_, shiftedA_4__22_, shiftedA_4__21_, 
        shiftedA_4__20_, shiftedA_4__19_, shiftedA_4__18_, shiftedA_4__17_, 
        shiftedA_4__16_, shiftedA_4__15_, shiftedA_4__14_, shiftedA_4__13_, 
        shiftedA_4__12_, shiftedA_4__11_, shiftedA_4__10_, shiftedA_4__9_, 
        shiftedA_4__8_, shiftedA_4__7_, shiftedA_4__6_, shiftedA_4__5_, 
        shiftedA_4__4_, 1'b0, 1'b0, 1'b0, 1'b0}), .c({n363, n363, n363, n363, 
        n362, n362, n362, n362, n362, n362, n362, n362, n362, n362, n362, n362, 
        n361, n361, n361, n361, n361, n361, n361, n361, n361, n361, n361, n361, 
        shiftedA_5__35_, shiftedA_5__34_, shiftedA_5__33_, shiftedA_5__32_, 
        shiftedA_5__31_, shiftedA_5__30_, shiftedA_5__29_, shiftedA_5__28_, 
        shiftedA_5__27_, shiftedA_5__26_, shiftedA_5__25_, shiftedA_5__24_, 
        shiftedA_5__23_, shiftedA_5__22_, shiftedA_5__21_, shiftedA_5__20_, 
        shiftedA_5__19_, shiftedA_5__18_, shiftedA_5__17_, shiftedA_5__16_, 
        shiftedA_5__15_, shiftedA_5__14_, shiftedA_5__13_, shiftedA_5__12_, 
        shiftedA_5__11_, shiftedA_5__10_, shiftedA_5__9_, shiftedA_5__8_, 
        shiftedA_5__7_, shiftedA_5__6_, shiftedA_5__5_, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .result(adderResult_level1[127:64]), .carry(
        carry_level1[127:64]) );
  BWAdder_60 level1_2__adder ( .a({n366, n366, n366, n365, n365, n365, n365, 
        n365, n365, n365, n365, n365, n365, n365, n365, n364, n364, n364, n364, 
        n364, n364, n364, n364, n364, n364, n364, n364, shiftedA_6__36_, 
        shiftedA_6__35_, shiftedA_6__34_, shiftedA_6__33_, shiftedA_6__32_, 
        shiftedA_6__31_, shiftedA_6__30_, shiftedA_6__29_, shiftedA_6__28_, 
        shiftedA_6__27_, shiftedA_6__26_, shiftedA_6__25_, shiftedA_6__24_, 
        shiftedA_6__23_, shiftedA_6__22_, shiftedA_6__21_, shiftedA_6__20_, 
        shiftedA_6__19_, shiftedA_6__18_, shiftedA_6__17_, shiftedA_6__16_, 
        shiftedA_6__15_, shiftedA_6__14_, shiftedA_6__13_, shiftedA_6__12_, 
        shiftedA_6__11_, shiftedA_6__10_, shiftedA_6__9_, shiftedA_6__8_, 
        shiftedA_6__7_, shiftedA_6__6_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .b({n369, n369, n368, n368, n368, n368, n368, n368, n368, n368, n368, 
        n368, n368, n368, n367, n367, n367, n367, n367, n367, n367, n367, n367, 
        n367, n367, n367, shiftedA_7__37_, shiftedA_7__36_, shiftedA_7__35_, 
        shiftedA_7__34_, shiftedA_7__33_, shiftedA_7__32_, shiftedA_7__31_, 
        shiftedA_7__30_, shiftedA_7__29_, shiftedA_7__28_, shiftedA_7__27_, 
        shiftedA_7__26_, shiftedA_7__25_, shiftedA_7__24_, shiftedA_7__23_, 
        shiftedA_7__22_, shiftedA_7__21_, shiftedA_7__20_, shiftedA_7__19_, 
        shiftedA_7__18_, shiftedA_7__17_, shiftedA_7__16_, shiftedA_7__15_, 
        shiftedA_7__14_, shiftedA_7__13_, shiftedA_7__12_, shiftedA_7__11_, 
        shiftedA_7__10_, shiftedA_7__9_, shiftedA_7__8_, shiftedA_7__7_, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({n259, n259, n259, n259, n259, 
        n259, n259, n258, n258, n258, n258, n258, n258, n257, n257, n257, n257, 
        n257, n257, n256, n256, n256, n256, n256, n256, shiftedA_8__38_, 
        shiftedA_8__37_, shiftedA_8__36_, shiftedA_8__35_, shiftedA_8__34_, 
        shiftedA_8__33_, shiftedA_8__32_, shiftedA_8__31_, shiftedA_8__30_, 
        shiftedA_8__29_, shiftedA_8__28_, shiftedA_8__27_, shiftedA_8__26_, 
        shiftedA_8__25_, shiftedA_8__24_, shiftedA_8__23_, shiftedA_8__22_, 
        shiftedA_8__21_, shiftedA_8__20_, shiftedA_8__19_, shiftedA_8__18_, 
        shiftedA_8__17_, shiftedA_8__16_, shiftedA_8__15_, shiftedA_8__14_, 
        shiftedA_8__13_, shiftedA_8__12_, shiftedA_8__11_, shiftedA_8__10_, 
        shiftedA_8__9_, shiftedA_8__8_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .result(adderResult_level1[191:128]), .carry(
        carry_level1[191:128]) );
  BWAdder_59 level1_3__adder ( .a({n261, n261, n261, n261, n261, n261, n261, 
        n261, n261, n261, n261, n261, n260, n260, n260, n260, n260, n260, n260, 
        n260, n260, n260, n260, n260, shiftedA_9__39_, shiftedA_9__38_, 
        shiftedA_9__37_, shiftedA_9__36_, shiftedA_9__35_, shiftedA_9__34_, 
        shiftedA_9__33_, shiftedA_9__32_, shiftedA_9__31_, shiftedA_9__30_, 
        shiftedA_9__29_, shiftedA_9__28_, shiftedA_9__27_, shiftedA_9__26_, 
        shiftedA_9__25_, shiftedA_9__24_, shiftedA_9__23_, shiftedA_9__22_, 
        shiftedA_9__21_, shiftedA_9__20_, shiftedA_9__19_, shiftedA_9__18_, 
        shiftedA_9__17_, shiftedA_9__16_, shiftedA_9__15_, shiftedA_9__14_, 
        shiftedA_9__13_, shiftedA_9__12_, shiftedA_9__11_, shiftedA_9__10_, 
        shiftedA_9__9_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .b({n263, n263, n263, n263, n263, n263, n263, n263, n263, n263, n263, 
        n262, n262, n262, n262, n262, n262, n262, n262, n262, n262, n262, n262, 
        shiftedA_10__40_, shiftedA_10__39_, shiftedA_10__38_, shiftedA_10__37_, 
        shiftedA_10__36_, shiftedA_10__35_, shiftedA_10__34_, shiftedA_10__33_, 
        shiftedA_10__32_, shiftedA_10__31_, shiftedA_10__30_, shiftedA_10__29_, 
        shiftedA_10__28_, shiftedA_10__27_, shiftedA_10__26_, shiftedA_10__25_, 
        shiftedA_10__24_, shiftedA_10__23_, shiftedA_10__22_, shiftedA_10__21_, 
        shiftedA_10__20_, shiftedA_10__19_, shiftedA_10__18_, shiftedA_10__17_, 
        shiftedA_10__16_, shiftedA_10__15_, shiftedA_10__14_, shiftedA_10__13_, 
        shiftedA_10__12_, shiftedA_10__11_, shiftedA_10__10_, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({n265, n265, n265, n265, 
        n265, n265, n265, n265, n265, n265, n264, n264, n264, n264, n264, n264, 
        n264, n264, n264, n264, n264, n264, shiftedA_11__41_, shiftedA_11__40_, 
        shiftedA_11__39_, shiftedA_11__38_, shiftedA_11__37_, shiftedA_11__36_, 
        shiftedA_11__35_, shiftedA_11__34_, shiftedA_11__33_, shiftedA_11__32_, 
        shiftedA_11__31_, shiftedA_11__30_, shiftedA_11__29_, shiftedA_11__28_, 
        shiftedA_11__27_, shiftedA_11__26_, shiftedA_11__25_, shiftedA_11__24_, 
        shiftedA_11__23_, shiftedA_11__22_, shiftedA_11__21_, shiftedA_11__20_, 
        shiftedA_11__19_, shiftedA_11__18_, shiftedA_11__17_, shiftedA_11__16_, 
        shiftedA_11__15_, shiftedA_11__14_, shiftedA_11__13_, shiftedA_11__12_, 
        shiftedA_11__11_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .result(adderResult_level1[255:192]), .carry(
        carry_level1[255:192]) );
  BWAdder_58 level1_4__adder ( .a({n267, n267, n267, n267, n267, n267, n267, 
        n267, n267, n266, n266, n266, n266, n266, n266, n266, n266, n266, n266, 
        n266, n266, shiftedA_12__42_, shiftedA_12__41_, shiftedA_12__40_, 
        shiftedA_12__39_, shiftedA_12__38_, shiftedA_12__37_, shiftedA_12__36_, 
        shiftedA_12__35_, shiftedA_12__34_, shiftedA_12__33_, shiftedA_12__32_, 
        shiftedA_12__31_, shiftedA_12__30_, shiftedA_12__29_, shiftedA_12__28_, 
        shiftedA_12__27_, shiftedA_12__26_, shiftedA_12__25_, shiftedA_12__24_, 
        shiftedA_12__23_, shiftedA_12__22_, shiftedA_12__21_, shiftedA_12__20_, 
        shiftedA_12__19_, shiftedA_12__18_, shiftedA_12__17_, shiftedA_12__16_, 
        shiftedA_12__15_, shiftedA_12__14_, shiftedA_12__13_, shiftedA_12__12_, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n269, n269, n269, n269, n269, n269, n269, n269, n268, n268, n268, n268, 
        n268, n268, n268, n268, n268, n268, n268, n268, shiftedA_13__43_, 
        shiftedA_13__42_, shiftedA_13__41_, shiftedA_13__40_, shiftedA_13__39_, 
        shiftedA_13__38_, shiftedA_13__37_, shiftedA_13__36_, shiftedA_13__35_, 
        shiftedA_13__34_, shiftedA_13__33_, shiftedA_13__32_, shiftedA_13__31_, 
        shiftedA_13__30_, shiftedA_13__29_, shiftedA_13__28_, shiftedA_13__27_, 
        shiftedA_13__26_, shiftedA_13__25_, shiftedA_13__24_, shiftedA_13__23_, 
        shiftedA_13__22_, shiftedA_13__21_, shiftedA_13__20_, shiftedA_13__19_, 
        shiftedA_13__18_, shiftedA_13__17_, shiftedA_13__16_, shiftedA_13__15_, 
        shiftedA_13__14_, shiftedA_13__13_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({n271, n271, n271, n271, 
        n271, n271, n271, n270, n270, n270, n270, n270, n270, n270, n270, n270, 
        n270, n270, n270, shiftedA_14__44_, shiftedA_14__43_, shiftedA_14__42_, 
        shiftedA_14__41_, shiftedA_14__40_, shiftedA_14__39_, shiftedA_14__38_, 
        shiftedA_14__37_, shiftedA_14__36_, shiftedA_14__35_, shiftedA_14__34_, 
        shiftedA_14__33_, shiftedA_14__32_, shiftedA_14__31_, shiftedA_14__30_, 
        shiftedA_14__29_, shiftedA_14__28_, shiftedA_14__27_, shiftedA_14__26_, 
        shiftedA_14__25_, shiftedA_14__24_, shiftedA_14__23_, shiftedA_14__22_, 
        shiftedA_14__21_, shiftedA_14__20_, shiftedA_14__19_, shiftedA_14__18_, 
        shiftedA_14__17_, shiftedA_14__16_, shiftedA_14__15_, shiftedA_14__14_, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .result(adderResult_level1[319:256]), .carry(
        carry_level1[319:256]) );
  BWAdder_57 level1_5__adder ( .a({n274, n274, n274, n274, n274, n274, n273, 
        n273, n273, n273, n273, n273, n272, n272, n272, n272, n272, n272, 
        shiftedA_15__45_, shiftedA_15__44_, shiftedA_15__43_, shiftedA_15__42_, 
        shiftedA_15__41_, shiftedA_15__40_, shiftedA_15__39_, shiftedA_15__38_, 
        shiftedA_15__37_, shiftedA_15__36_, shiftedA_15__35_, shiftedA_15__34_, 
        shiftedA_15__33_, shiftedA_15__32_, shiftedA_15__31_, shiftedA_15__30_, 
        shiftedA_15__29_, shiftedA_15__28_, shiftedA_15__27_, shiftedA_15__26_, 
        shiftedA_15__25_, shiftedA_15__24_, shiftedA_15__23_, shiftedA_15__22_, 
        shiftedA_15__21_, shiftedA_15__20_, shiftedA_15__19_, shiftedA_15__18_, 
        shiftedA_15__17_, shiftedA_15__16_, shiftedA_15__15_, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n277, n277, n277, n277, n277, n276, n276, n276, n276, n276, n276, n275, 
        n275, n275, n275, n275, n275, shiftedA_16__46_, shiftedA_16__45_, 
        shiftedA_16__44_, shiftedA_16__43_, shiftedA_16__42_, shiftedA_16__41_, 
        shiftedA_16__40_, shiftedA_16__39_, shiftedA_16__38_, shiftedA_16__37_, 
        shiftedA_16__36_, shiftedA_16__35_, shiftedA_16__34_, shiftedA_16__33_, 
        shiftedA_16__32_, shiftedA_16__31_, shiftedA_16__30_, shiftedA_16__29_, 
        shiftedA_16__28_, shiftedA_16__27_, shiftedA_16__26_, shiftedA_16__25_, 
        shiftedA_16__24_, shiftedA_16__23_, shiftedA_16__22_, shiftedA_16__21_, 
        shiftedA_16__20_, shiftedA_16__19_, shiftedA_16__18_, shiftedA_16__17_, 
        shiftedA_16__16_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({n280, n280, n280, n280, 
        n279, n279, n279, n279, n279, n279, n278, n278, n278, n278, n278, n278, 
        shiftedA_17__47_, shiftedA_17__46_, shiftedA_17__45_, shiftedA_17__44_, 
        shiftedA_17__43_, shiftedA_17__42_, shiftedA_17__41_, shiftedA_17__40_, 
        shiftedA_17__39_, shiftedA_17__38_, shiftedA_17__37_, shiftedA_17__36_, 
        shiftedA_17__35_, shiftedA_17__34_, shiftedA_17__33_, shiftedA_17__32_, 
        shiftedA_17__31_, shiftedA_17__30_, shiftedA_17__29_, shiftedA_17__28_, 
        shiftedA_17__27_, shiftedA_17__26_, shiftedA_17__25_, shiftedA_17__24_, 
        shiftedA_17__23_, shiftedA_17__22_, shiftedA_17__21_, shiftedA_17__20_, 
        shiftedA_17__19_, shiftedA_17__18_, shiftedA_17__17_, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .result(adderResult_level1[383:320]), .carry(
        carry_level1[383:320]) );
  BWAdder_56 level1_6__adder ( .a({n283, n283, n283, n282, n282, n282, n282, 
        n282, n282, n281, n281, n281, n281, n281, n281, shiftedA_18__48_, 
        shiftedA_18__47_, shiftedA_18__46_, shiftedA_18__45_, shiftedA_18__44_, 
        shiftedA_18__43_, shiftedA_18__42_, shiftedA_18__41_, shiftedA_18__40_, 
        shiftedA_18__39_, shiftedA_18__38_, shiftedA_18__37_, shiftedA_18__36_, 
        shiftedA_18__35_, shiftedA_18__34_, shiftedA_18__33_, shiftedA_18__32_, 
        shiftedA_18__31_, shiftedA_18__30_, shiftedA_18__29_, shiftedA_18__28_, 
        shiftedA_18__27_, shiftedA_18__26_, shiftedA_18__25_, shiftedA_18__24_, 
        shiftedA_18__23_, shiftedA_18__22_, shiftedA_18__21_, shiftedA_18__20_, 
        shiftedA_18__19_, shiftedA_18__18_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n286, n286, n285, n285, n285, n285, n285, n285, n284, n284, n284, n284, 
        n284, n284, shiftedA_19__49_, shiftedA_19__48_, shiftedA_19__47_, 
        shiftedA_19__46_, shiftedA_19__45_, shiftedA_19__44_, shiftedA_19__43_, 
        shiftedA_19__42_, shiftedA_19__41_, shiftedA_19__40_, shiftedA_19__39_, 
        shiftedA_19__38_, shiftedA_19__37_, shiftedA_19__36_, shiftedA_19__35_, 
        shiftedA_19__34_, shiftedA_19__33_, shiftedA_19__32_, shiftedA_19__31_, 
        shiftedA_19__30_, shiftedA_19__29_, shiftedA_19__28_, shiftedA_19__27_, 
        shiftedA_19__26_, shiftedA_19__25_, shiftedA_19__24_, shiftedA_19__23_, 
        shiftedA_19__22_, shiftedA_19__21_, shiftedA_19__20_, shiftedA_19__19_, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({n288, n288, n288, n288, 
        n288, n288, n288, n287, n287, n287, n287, n287, n287, shiftedA_20__50_, 
        shiftedA_20__49_, shiftedA_20__48_, shiftedA_20__47_, shiftedA_20__46_, 
        shiftedA_20__45_, shiftedA_20__44_, shiftedA_20__43_, shiftedA_20__42_, 
        shiftedA_20__41_, shiftedA_20__40_, shiftedA_20__39_, shiftedA_20__38_, 
        shiftedA_20__37_, shiftedA_20__36_, shiftedA_20__35_, shiftedA_20__34_, 
        shiftedA_20__33_, shiftedA_20__32_, shiftedA_20__31_, shiftedA_20__30_, 
        shiftedA_20__29_, shiftedA_20__28_, shiftedA_20__27_, shiftedA_20__26_, 
        shiftedA_20__25_, shiftedA_20__24_, shiftedA_20__23_, shiftedA_20__22_, 
        shiftedA_20__21_, shiftedA_20__20_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .result(adderResult_level1[447:384]), .carry(
        carry_level1[447:384]) );
  BWAdder_55 level1_7__adder ( .a({shiftedA_21__63_, shiftedA_21__63_, 
        shiftedA_21__63_, shiftedA_21__63_, shiftedA_21__63_, shiftedA_21__63_, 
        shiftedA_21__63_, shiftedA_21__63_, shiftedA_21__63_, shiftedA_21__63_, 
        shiftedA_21__63_, shiftedA_21__63_, shiftedA_21__51_, shiftedA_21__50_, 
        shiftedA_21__49_, shiftedA_21__48_, shiftedA_21__47_, shiftedA_21__46_, 
        shiftedA_21__45_, shiftedA_21__44_, shiftedA_21__43_, shiftedA_21__42_, 
        shiftedA_21__41_, shiftedA_21__40_, shiftedA_21__39_, shiftedA_21__38_, 
        shiftedA_21__37_, shiftedA_21__36_, shiftedA_21__35_, shiftedA_21__34_, 
        shiftedA_21__33_, shiftedA_21__32_, shiftedA_21__31_, shiftedA_21__30_, 
        shiftedA_21__29_, shiftedA_21__28_, shiftedA_21__27_, shiftedA_21__26_, 
        shiftedA_21__25_, shiftedA_21__24_, shiftedA_21__23_, shiftedA_21__22_, 
        shiftedA_21__21_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_22__63_, shiftedA_22__63_, shiftedA_22__63_, shiftedA_22__63_, 
        shiftedA_22__63_, shiftedA_22__63_, shiftedA_22__63_, shiftedA_22__63_, 
        shiftedA_22__63_, shiftedA_22__63_, shiftedA_22__63_, shiftedA_22__52_, 
        shiftedA_22__51_, shiftedA_22__50_, shiftedA_22__49_, shiftedA_22__48_, 
        shiftedA_22__47_, shiftedA_22__46_, shiftedA_22__45_, shiftedA_22__44_, 
        shiftedA_22__43_, shiftedA_22__42_, shiftedA_22__41_, shiftedA_22__40_, 
        shiftedA_22__39_, shiftedA_22__38_, shiftedA_22__37_, shiftedA_22__36_, 
        shiftedA_22__35_, shiftedA_22__34_, shiftedA_22__33_, shiftedA_22__32_, 
        shiftedA_22__31_, shiftedA_22__30_, shiftedA_22__29_, shiftedA_22__28_, 
        shiftedA_22__27_, shiftedA_22__26_, shiftedA_22__25_, shiftedA_22__24_, 
        shiftedA_22__23_, shiftedA_22__22_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_23__63_, shiftedA_23__63_, 
        shiftedA_23__63_, shiftedA_23__63_, shiftedA_23__63_, shiftedA_23__63_, 
        shiftedA_23__63_, shiftedA_23__63_, shiftedA_23__63_, shiftedA_23__63_, 
        shiftedA_23__53_, shiftedA_23__52_, shiftedA_23__51_, shiftedA_23__50_, 
        shiftedA_23__49_, shiftedA_23__48_, shiftedA_23__47_, shiftedA_23__46_, 
        shiftedA_23__45_, shiftedA_23__44_, shiftedA_23__43_, shiftedA_23__42_, 
        shiftedA_23__41_, shiftedA_23__40_, shiftedA_23__39_, shiftedA_23__38_, 
        shiftedA_23__37_, shiftedA_23__36_, shiftedA_23__35_, shiftedA_23__34_, 
        shiftedA_23__33_, shiftedA_23__32_, shiftedA_23__31_, shiftedA_23__30_, 
        shiftedA_23__29_, shiftedA_23__28_, shiftedA_23__27_, shiftedA_23__26_, 
        shiftedA_23__25_, shiftedA_23__24_, shiftedA_23__23_, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[511:448]), .carry(carry_level1[511:448]) );
  BWAdder_54 level1_8__adder ( .a({shiftedA_24__63_, shiftedA_24__63_, 
        shiftedA_24__63_, shiftedA_24__63_, shiftedA_24__63_, shiftedA_24__63_, 
        shiftedA_24__63_, shiftedA_24__63_, shiftedA_24__63_, shiftedA_24__54_, 
        shiftedA_24__53_, shiftedA_24__52_, shiftedA_24__51_, shiftedA_24__50_, 
        shiftedA_24__49_, shiftedA_24__48_, shiftedA_24__47_, shiftedA_24__46_, 
        shiftedA_24__45_, shiftedA_24__44_, shiftedA_24__43_, shiftedA_24__42_, 
        shiftedA_24__41_, shiftedA_24__40_, shiftedA_24__39_, shiftedA_24__38_, 
        shiftedA_24__37_, shiftedA_24__36_, shiftedA_24__35_, shiftedA_24__34_, 
        shiftedA_24__33_, shiftedA_24__32_, shiftedA_24__31_, shiftedA_24__30_, 
        shiftedA_24__29_, shiftedA_24__28_, shiftedA_24__27_, shiftedA_24__26_, 
        shiftedA_24__25_, shiftedA_24__24_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_25__63_, 
        shiftedA_25__63_, shiftedA_25__63_, shiftedA_25__63_, shiftedA_25__63_, 
        shiftedA_25__63_, shiftedA_25__63_, shiftedA_25__63_, shiftedA_25__55_, 
        shiftedA_25__54_, shiftedA_25__53_, shiftedA_25__52_, shiftedA_25__51_, 
        shiftedA_25__50_, shiftedA_25__49_, shiftedA_25__48_, shiftedA_25__47_, 
        shiftedA_25__46_, shiftedA_25__45_, shiftedA_25__44_, shiftedA_25__43_, 
        shiftedA_25__42_, shiftedA_25__41_, shiftedA_25__40_, shiftedA_25__39_, 
        shiftedA_25__38_, shiftedA_25__37_, shiftedA_25__36_, shiftedA_25__35_, 
        shiftedA_25__34_, shiftedA_25__33_, shiftedA_25__32_, shiftedA_25__31_, 
        shiftedA_25__30_, shiftedA_25__29_, shiftedA_25__28_, shiftedA_25__27_, 
        shiftedA_25__26_, shiftedA_25__25_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_26__63_, 
        shiftedA_26__63_, shiftedA_26__63_, shiftedA_26__63_, shiftedA_26__63_, 
        shiftedA_26__63_, shiftedA_26__63_, shiftedA_26__56_, shiftedA_26__55_, 
        shiftedA_26__54_, shiftedA_26__53_, shiftedA_26__52_, shiftedA_26__51_, 
        shiftedA_26__50_, shiftedA_26__49_, shiftedA_26__48_, shiftedA_26__47_, 
        shiftedA_26__46_, shiftedA_26__45_, shiftedA_26__44_, shiftedA_26__43_, 
        shiftedA_26__42_, shiftedA_26__41_, shiftedA_26__40_, shiftedA_26__39_, 
        shiftedA_26__38_, shiftedA_26__37_, shiftedA_26__36_, shiftedA_26__35_, 
        shiftedA_26__34_, shiftedA_26__33_, shiftedA_26__32_, shiftedA_26__31_, 
        shiftedA_26__30_, shiftedA_26__29_, shiftedA_26__28_, shiftedA_26__27_, 
        shiftedA_26__26_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(adderResult_level1[575:512]), 
        .carry(carry_level1[575:512]) );
  BWAdder_53 level1_9__adder ( .a({shiftedA_27__63_, shiftedA_27__63_, 
        shiftedA_27__63_, shiftedA_27__63_, shiftedA_27__63_, shiftedA_27__63_, 
        shiftedA_27__57_, shiftedA_27__56_, shiftedA_27__55_, shiftedA_27__54_, 
        shiftedA_27__53_, shiftedA_27__52_, shiftedA_27__51_, shiftedA_27__50_, 
        shiftedA_27__49_, shiftedA_27__48_, shiftedA_27__47_, shiftedA_27__46_, 
        shiftedA_27__45_, shiftedA_27__44_, shiftedA_27__43_, shiftedA_27__42_, 
        shiftedA_27__41_, shiftedA_27__40_, shiftedA_27__39_, shiftedA_27__38_, 
        shiftedA_27__37_, shiftedA_27__36_, shiftedA_27__35_, shiftedA_27__34_, 
        shiftedA_27__33_, shiftedA_27__32_, shiftedA_27__31_, shiftedA_27__30_, 
        shiftedA_27__29_, shiftedA_27__28_, shiftedA_27__27_, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_28__63_, shiftedA_28__63_, shiftedA_28__63_, shiftedA_28__63_, 
        shiftedA_28__63_, shiftedA_28__58_, shiftedA_28__57_, shiftedA_28__56_, 
        shiftedA_28__55_, shiftedA_28__54_, shiftedA_28__53_, shiftedA_28__52_, 
        shiftedA_28__51_, shiftedA_28__50_, shiftedA_28__49_, shiftedA_28__48_, 
        shiftedA_28__47_, shiftedA_28__46_, shiftedA_28__45_, shiftedA_28__44_, 
        shiftedA_28__43_, shiftedA_28__42_, shiftedA_28__41_, shiftedA_28__40_, 
        shiftedA_28__39_, shiftedA_28__38_, shiftedA_28__37_, shiftedA_28__36_, 
        shiftedA_28__35_, shiftedA_28__34_, shiftedA_28__33_, shiftedA_28__32_, 
        shiftedA_28__31_, shiftedA_28__30_, shiftedA_28__29_, shiftedA_28__28_, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_29__63_, shiftedA_29__63_, 
        shiftedA_29__63_, shiftedA_29__63_, shiftedA_29__59_, shiftedA_29__58_, 
        shiftedA_29__57_, shiftedA_29__56_, shiftedA_29__55_, shiftedA_29__54_, 
        shiftedA_29__53_, shiftedA_29__52_, shiftedA_29__51_, shiftedA_29__50_, 
        shiftedA_29__49_, shiftedA_29__48_, shiftedA_29__47_, shiftedA_29__46_, 
        shiftedA_29__45_, shiftedA_29__44_, shiftedA_29__43_, shiftedA_29__42_, 
        shiftedA_29__41_, shiftedA_29__40_, shiftedA_29__39_, shiftedA_29__38_, 
        shiftedA_29__37_, shiftedA_29__36_, shiftedA_29__35_, shiftedA_29__34_, 
        shiftedA_29__33_, shiftedA_29__32_, shiftedA_29__31_, shiftedA_29__30_, 
        shiftedA_29__29_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[639:576]), .carry(carry_level1[639:576]) );
  BWAdder_52 level1_10__adder ( .a({shiftedA_30__63_, shiftedA_30__63_, 
        shiftedA_30__63_, shiftedA_30__60_, shiftedA_30__59_, shiftedA_30__58_, 
        shiftedA_30__57_, shiftedA_30__56_, shiftedA_30__55_, shiftedA_30__54_, 
        shiftedA_30__53_, shiftedA_30__52_, shiftedA_30__51_, shiftedA_30__50_, 
        shiftedA_30__49_, shiftedA_30__48_, shiftedA_30__47_, shiftedA_30__46_, 
        shiftedA_30__45_, shiftedA_30__44_, shiftedA_30__43_, shiftedA_30__42_, 
        shiftedA_30__41_, shiftedA_30__40_, shiftedA_30__39_, shiftedA_30__38_, 
        shiftedA_30__37_, shiftedA_30__36_, shiftedA_30__35_, shiftedA_30__34_, 
        shiftedA_30__33_, shiftedA_30__32_, shiftedA_30__31_, shiftedA_30__30_, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_32__63_, 
        shiftedA_32__63_, shiftedA_33__63_, shiftedA_34__63_, shiftedA_35__63_, 
        shiftedA_36__63_, shiftedA_37__63_, shiftedA_38__63_, shiftedA_39__63_, 
        shiftedA_40__63_, shiftedA_41__63_, shiftedA_42__63_, n290, n292, n296, 
        n299, n302, n305, n307, n309, n311, n313, n315, n317, n320, n323, n327, 
        n329, n333, n336, n338, n342, n345, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .c({shiftedA_32__63_, shiftedA_33__63_, shiftedA_34__63_, 
        shiftedA_35__63_, shiftedA_36__63_, shiftedA_37__63_, shiftedA_38__63_, 
        shiftedA_39__63_, shiftedA_40__63_, shiftedA_41__63_, shiftedA_42__63_, 
        n289, n291, n294, n297, n300, n303, n306, n308, n310, n312, n314, n316, 
        n318, n322, n325, n328, n331, n334, n337, n340, n343, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(adderResult_level1[703:640]), 
        .carry(carry_level1[703:640]) );
  BWAdder_51 level1_11__adder ( .a({shiftedA_33__63_, shiftedA_34__63_, 
        shiftedA_35__63_, shiftedA_36__63_, shiftedA_37__63_, shiftedA_38__63_, 
        shiftedA_39__63_, shiftedA_40__63_, shiftedA_41__63_, shiftedA_42__63_, 
        n289, n291, n294, n298, n301, n304, n306, n308, n311, n313, n315, n316, 
        n319, n322, n326, n328, n332, n335, n337, n341, n344, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_34__63_, 
        shiftedA_35__63_, shiftedA_36__63_, shiftedA_37__63_, shiftedA_38__63_, 
        shiftedA_39__63_, shiftedA_40__63_, shiftedA_41__63_, shiftedA_42__63_, 
        n290, n292, n296, n299, n302, n305, n307, n309, n311, n313, n315, n317, 
        n321, n323, n327, n330, n333, n336, n339, n342, n345, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_35__63_, 
        shiftedA_36__63_, shiftedA_37__63_, shiftedA_38__63_, shiftedA_39__63_, 
        shiftedA_40__63_, shiftedA_41__63_, shiftedA_42__63_, n289, n291, n294, 
        n297, n300, n303, n306, n308, n310, n312, n314, n316, n318, n322, n325, 
        n328, n331, n334, n337, n340, n343, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(adderResult_level1[767:704]), 
        .carry(carry_level1[767:704]) );
  BWAdder_50 level1_12__adder ( .a({shiftedA_36__63_, shiftedA_37__63_, 
        shiftedA_38__63_, shiftedA_39__63_, shiftedA_40__63_, shiftedA_41__63_, 
        shiftedA_42__63_, n290, n292, n295, n297, n301, n304, n306, n308, n310, 
        n313, n315, n316, n319, n322, n326, n328, n332, n334, n338, n341, n344, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_37__63_, shiftedA_38__63_, shiftedA_39__63_, shiftedA_40__63_, 
        shiftedA_41__63_, shiftedA_42__63_, n290, n292, n295, n298, n301, n305, 
        n307, n309, n311, n313, n315, n317, n321, n323, n326, n330, n332, n335, 
        n339, n342, n345, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_38__63_, shiftedA_39__63_, 
        shiftedA_40__63_, shiftedA_41__63_, shiftedA_42__63_, n289, n291, n294, 
        n297, n300, n303, n306, n308, n310, n312, n314, n316, n318, n322, n325, 
        n328, n331, n334, n337, n340, n343, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[831:768]), .carry(carry_level1[831:768]) );
  BWAdder_49 level1_13__adder ( .a({shiftedA_39__63_, shiftedA_40__63_, 
        shiftedA_41__63_, shiftedA_42__63_, n290, n292, n295, n298, n301, n304, 
        n306, n308, n310, n312, n314, n316, n320, n323, n326, n328, n332, n334, 
        n338, n341, n344, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_40__63_, 
        shiftedA_41__63_, shiftedA_42__63_, n290, n292, n295, n298, n301, n304, 
        n307, n309, n311, n313, n315, n317, n321, n324, n326, n330, n332, n335, 
        n339, n342, n345, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_41__63_, 
        shiftedA_42__63_, n289, n291, n294, n297, n300, n303, n306, n308, n310, 
        n312, n314, n316, n318, n322, n325, n328, n331, n334, n337, n340, n343, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(adderResult_level1[895:832]), 
        .carry(carry_level1[895:832]) );
  BWAdder_48 level1_14__adder ( .a({shiftedA_42__63_, n289, n291, n295, n298, 
        n301, n304, n306, n308, n310, n312, n314, n316, n320, n323, n326, n329, 
        n332, n335, n338, n341, n344, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .b({n289, n293, n295, n299, n302, n305, n307, n309, n311, n313, n315, 
        n317, n321, n323, n326, n329, n332, n335, n339, n341, n345, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({n293, n294, n297, n300, n303, n306, 
        n308, n310, n312, n314, n316, n319, n322, n325, n328, n331, n334, n337, 
        n340, n343, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[959:896]), .carry(carry_level1[959:896]) );
  BWAdder_47 level1_15__adder ( .a({n296, n298, n300, n304, n306, n308, n310, 
        n312, n314, n317, n320, n323, n325, n329, n331, n335, n338, n341, n344, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n299, n302, 
        n305, n307, n309, n311, n313, n315, n317, n321, n323, n326, n329, n332, 
        n335, n339, n341, n344, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .c({n302, n303, n306, n308, n310, n312, n314, n316, n319, 
        n322, n325, n328, n331, n334, n337, n340, n343, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[1023:960]), .carry(carry_level1[1023:960]) );
  BWAdder_46 level1_16__adder ( .a({n305, n306, n308, n310, n312, n314, n317, 
        n319, n323, n326, n329, n332, n335, n338, n341, n344, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n307, n309, 
        n311, n313, n315, n317, n321, n323, n326, n329, n332, n335, n339, n341, 
        n344, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .c({n309, n310, n312, n314, n316, n318, n322, n325, n328, 
        n331, n334, n337, n340, n343, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[1087:1024]), .carry(carry_level1[1087:1024]) );
  BWAdder_45 level1_17__adder ( .a({n311, n312, n314, n317, n319, n322, n325, 
        n329, n331, n335, n338, n340, n344, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n313, n315, 
        n317, n320, n323, n326, n329, n332, n336, n338, n341, n344, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .c({n315, n316, n318, n322, n325, n328, n331, n334, n337, 
        n340, n343, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[1151:1088]), .carry(carry_level1[1151:1088]) );
  BWAdder_44 level1_18__adder ( .a({n317, n320, n322, n325, n329, n331, n335, 
        n338, n341, n344, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n321, n323, 
        n326, n329, n333, n336, n338, n342, n345, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .c({n324, n325, n328, n331, n334, n337, n340, n343, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[1215:1152]), .carry(carry_level1[1215:1152]) );
  BWAdder_43 level1_19__adder ( .a({n327, n329, n332, n335, n337, n340, n343, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n330, n333, 
        n336, n338, n342, n345, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .c({n333, n334, n337, n340, n343, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[1279:1216]), .carry(carry_level1[1279:1216]) );
  BWAdder_42 level1_20__adder ( .a({n336, n338, n341, n344, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n339, n342, 
        n345, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .c({n342, n343, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[1343:1280]), .carry(carry_level1[1343:1280]) );
  BWAdder_41 level2_a_0__adder ( .a(adderResult_level1[63:0]), .b(
        adderResult_level1[127:64]), .c(adderResult_level1[191:128]), .result(
        adderResult_level2[63:0]), .carry(carry_level2[63:0]) );
  BWAdder_40 level2_a_1__adder ( .a(adderResult_level1[255:192]), .b(
        adderResult_level1[319:256]), .c(adderResult_level1[383:320]), 
        .result(adderResult_level2[127:64]), .carry(carry_level2[127:64]) );
  BWAdder_39 level2_a_2__adder ( .a(adderResult_level1[447:384]), .b(
        adderResult_level1[511:448]), .c(adderResult_level1[575:512]), 
        .result(adderResult_level2[191:128]), .carry(carry_level2[191:128]) );
  BWAdder_38 level2_a_3__adder ( .a(adderResult_level1[639:576]), .b(
        adderResult_level1[703:640]), .c(adderResult_level1[767:704]), 
        .result(adderResult_level2[255:192]), .carry(carry_level2[255:192]) );
  BWAdder_37 level2_a_4__adder ( .a(adderResult_level1[831:768]), .b(
        adderResult_level1[895:832]), .c(adderResult_level1[959:896]), 
        .result(adderResult_level2[319:256]), .carry(carry_level2[319:256]) );
  BWAdder_36 level2_a_5__adder ( .a(adderResult_level1[1023:960]), .b(
        adderResult_level1[1087:1024]), .c(adderResult_level1[1151:1088]), 
        .result(adderResult_level2[383:320]), .carry(carry_level2[383:320]) );
  BWAdder_35 level2_a_6__adder ( .a(adderResult_level1[1215:1152]), .b(
        adderResult_level1[1279:1216]), .c(adderResult_level1[1343:1280]), 
        .result(adderResult_level2[447:384]), .carry(carry_level2[447:384]) );
  BWAdder_34 level2_b_0__adder ( .a({carry_level1[63:1], 1'b0}), .b({
        carry_level1[127:65], 1'b0}), .c({carry_level1[191:129], 1'b0}), 
        .result(adderResult_level2[511:448]), .carry(carry_level2[511:448]) );
  BWAdder_33 level2_b_1__adder ( .a({carry_level1[255:193], 1'b0}), .b({
        carry_level1[319:257], 1'b0}), .c({carry_level1[383:321], 1'b0}), 
        .result(adderResult_level2[575:512]), .carry(carry_level2[575:512]) );
  BWAdder_32 level2_b_2__adder ( .a({carry_level1[447:385], 1'b0}), .b({
        carry_level1[511:449], 1'b0}), .c({carry_level1[575:513], 1'b0}), 
        .result(adderResult_level2[639:576]), .carry(carry_level2[639:576]) );
  BWAdder_31 level2_b_3__adder ( .a({carry_level1[639:577], 1'b0}), .b({
        carry_level1[703:641], 1'b0}), .c({carry_level1[767:705], 1'b0}), 
        .result(adderResult_level2[703:640]), .carry(carry_level2[703:640]) );
  BWAdder_30 level2_b_4__adder ( .a({carry_level1[831:769], 1'b0}), .b({
        carry_level1[895:833], 1'b0}), .c({carry_level1[959:897], 1'b0}), 
        .result(adderResult_level2[767:704]), .carry(carry_level2[767:704]) );
  BWAdder_29 level2_b_5__adder ( .a({carry_level1[1023:961], 1'b0}), .b({
        carry_level1[1087:1025], 1'b0}), .c({carry_level1[1151:1089], 1'b0}), 
        .result(adderResult_level2[831:768]), .carry(carry_level2[831:768]) );
  BWAdder_28 level2_b_6__adder ( .a({carry_level1[1215:1153], 1'b0}), .b({
        carry_level1[1279:1217], 1'b0}), .c({carry_level1[1343:1281], 1'b0}), 
        .result(adderResult_level2[895:832]), .carry(carry_level2[895:832]) );
  BWAdder_27 level3_a_0__adder ( .a(adderResult_level2[63:0]), .b(
        adderResult_level2[127:64]), .c(adderResult_level2[191:128]), .result(
        adderResult_level3[63:0]), .carry(carry_level3[63:0]) );
  BWAdder_26 level3_a_1__adder ( .a(adderResult_level2[255:192]), .b(
        adderResult_level2[319:256]), .c(adderResult_level2[383:320]), 
        .result(adderResult_level3[127:64]), .carry(carry_level3[127:64]) );
  BWAdder_25 level3_a_2__adder ( .a(adderResult_level2[447:384]), .b(
        adderResult_level2[511:448]), .c(adderResult_level2[575:512]), 
        .result(adderResult_level3[191:128]), .carry(carry_level3[191:128]) );
  BWAdder_24 level3_a_3__adder ( .a(adderResult_level2[639:576]), .b(
        adderResult_level2[703:640]), .c(adderResult_level2[767:704]), 
        .result(adderResult_level3[255:192]), .carry(carry_level3[255:192]) );
  BWAdder_23 level3_b_0__adder ( .a({carry_level2[63:1], 1'b0}), .b({
        carry_level2[127:65], 1'b0}), .c({carry_level2[191:129], 1'b0}), 
        .result(adderResult_level3[319:256]), .carry(carry_level3[319:256]) );
  BWAdder_22 level3_b_1__adder ( .a({carry_level2[255:193], 1'b0}), .b({
        carry_level2[319:257], 1'b0}), .c({carry_level2[383:321], 1'b0}), 
        .result(adderResult_level3[383:320]), .carry(carry_level3[383:320]) );
  BWAdder_21 level3_b_2__adder ( .a({carry_level2[447:385], 1'b0}), .b({
        carry_level2[511:449], 1'b0}), .c({carry_level2[575:513], 1'b0}), 
        .result(adderResult_level3[447:384]), .carry(carry_level3[447:384]) );
  BWAdder_20 level3_b_3__adder ( .a({carry_level2[639:577], 1'b0}), .b({
        carry_level2[703:641], 1'b0}), .c({carry_level2[767:705], 1'b0}), 
        .result(adderResult_level3[511:448]), .carry(carry_level3[511:448]) );
  BWAdder_19 adder ( .a(adderResult_level2[831:768]), .b(
        adderResult_level2[895:832]), .c({carry_level2[831:769], 1'b0}), 
        .result(adderResult_level3[575:512]), .carry(carry_level3[575:512]) );
  BWAdder_18 level4_a_0__adder ( .a(adderResult_level3[63:0]), .b(
        adderResult_level3[127:64]), .c(adderResult_level3[191:128]), .result(
        adderResult_level4[63:0]), .carry(carry_level4[63:0]) );
  BWAdder_17 level4_a_1__adder ( .a(adderResult_level3[255:192]), .b(
        adderResult_level3[319:256]), .c(adderResult_level3[383:320]), 
        .result(adderResult_level4[127:64]), .carry(carry_level4[127:64]) );
  BWAdder_16 level4_a_2__adder ( .a(adderResult_level3[447:384]), .b(
        adderResult_level3[511:448]), .c(adderResult_level3[575:512]), 
        .result(adderResult_level4[191:128]), .carry(carry_level4[191:128]) );
  BWAdder_15 level4_b_0__adder ( .a({carry_level3[63:1], 1'b0}), .b({
        carry_level3[127:65], 1'b0}), .c({carry_level3[191:129], 1'b0}), 
        .result(adderResult_level4[255:192]), .carry(carry_level4[255:192]) );
  BWAdder_14 level4_b_1__adder ( .a({carry_level3[255:193], 1'b0}), .b({
        carry_level3[319:257], 1'b0}), .c({carry_level3[383:321], 1'b0}), 
        .result(adderResult_level4[319:256]), .carry(carry_level4[319:256]) );
  BWAdder_13 level4_b_2__adder ( .a({carry_level3[447:385], 1'b0}), .b({
        carry_level3[511:449], 1'b0}), .c({carry_level3[575:513], 1'b0}), 
        .result(adderResult_level4[383:320]), .carry(carry_level4[383:320]) );
  BWAdder_12 level5_a_0__adder ( .a(adderResult_level4[63:0]), .b(
        adderResult_level4[127:64]), .c(adderResult_level4[191:128]), .result(
        adderResult_level5[63:0]), .carry(carry_level5[63:0]) );
  BWAdder_11 level5_a_1__adder ( .a(adderResult_level4[255:192]), .b(
        adderResult_level4[319:256]), .c(adderResult_level4[383:320]), 
        .result(adderResult_level5[127:64]), .carry(carry_level5[127:64]) );
  BWAdder_10 level5_b_0__adder ( .a({carry_level4[63:1], 1'b0}), .b({
        carry_level4[127:65], 1'b0}), .c({carry_level4[191:129], 1'b0}), 
        .result(adderResult_level5[191:128]), .carry(carry_level5[191:128]) );
  BWAdder_9 level5_b_1__adder ( .a({carry_level4[255:193], 1'b0}), .b({
        carry_level4[319:257], 1'b0}), .c({carry_level4[383:321], 1'b0}), 
        .result(adderResult_level5[255:192]), .carry(carry_level5[255:192]) );
  BWAdder_8 adder_0 ( .a(adderResult_level5[63:0]), .b(
        adderResult_level5[127:64]), .c(adderResult_level5[191:128]), .result(
        adderResult_level6[63:0]), .carry(carry_level6[63:0]) );
  BWAdder_7 adder_1 ( .a(adderResult_level5[255:192]), .b({carry_level5[63:1], 
        1'b0}), .c({carry_level5[127:65], 1'b0}), .result(
        adderResult_level6[127:64]), .carry(carry_level6[127:64]) );
  BWAdder_6 adder_2 ( .a({carry_level5[191:129], 1'b0}), .b({
        carry_level5[255:193], 1'b0}), .c({carry_level2[895:833], 1'b0}), 
        .result(adderResult_level6[191:128]), .carry(carry_level6[191:128]) );
  BWAdder_5 adder_3 ( .a(adderResult_level6[63:0]), .b(
        adderResult_level6[127:64]), .c(adderResult_level6[191:128]), .result(
        adderResult_level7[63:0]), .carry(carry_level7[63:0]) );
  BWAdder_4 adder_4 ( .a({carry_level6[63:1], 1'b0}), .b({carry_level6[127:65], 
        1'b0}), .c({carry_level6[191:129], 1'b0}), .result(
        adderResult_level7[127:64]), .carry(carry_level7[127:64]) );
  BWAdder_3 adder_5 ( .a(adderResult_level7[63:0]), .b(
        adderResult_level7[127:64]), .c({carry_level7[63:1], 1'b0}), .result(
        adderResult_level8), .carry(carry_level8) );
  BWAdder_2 adder_6 ( .a(adderResult_level8), .b({carry_level7[127:65], 1'b0}), 
        .c({carry_level8[63:1], 1'b0}), .result(adderResult_level9), .carry(
        carry_level9) );
  BWAdder_1 adder_7 ( .a(adderResult_level9), .b({n345, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .c({carry_level9[63:1], 1'b0}), .result(adderResult_level10), .carry(
        carry_level10) );
  CRAdder_64 CRAdd ( .a(adderResult_level10), .b({carry_level10[63:1], 1'b0}), 
        .cin(1'b0), .sum(result) );
  BUF_X4 U3 ( .A(n67), .Z(n80) );
  BUF_X1 U4 ( .A(n23), .Z(n189) );
  BUF_X2 U5 ( .A(n27), .Z(n179) );
  NOR2_X1 U6 ( .A1(n188), .A2(n86), .ZN(shiftedA_2__10_) );
  AND2_X1 U7 ( .A1(a[7]), .A2(n71), .ZN(shiftedA_0__7_) );
  BUF_X1 U8 ( .A(n61), .Z(n83) );
  AND2_X1 U9 ( .A1(b[22]), .A2(n374), .ZN(shiftedA_22__63_) );
  CLKBUF_X1 U10 ( .A(n63), .Z(n26) );
  BUF_X2 U11 ( .A(n61), .Z(n82) );
  CLKBUF_X1 U12 ( .A(n175), .Z(n29) );
  BUF_X2 U13 ( .A(n175), .Z(n63) );
  BUF_X1 U14 ( .A(n72), .Z(n175) );
  BUF_X2 U15 ( .A(n25), .Z(n183) );
  BUF_X2 U16 ( .A(n183), .Z(n182) );
  BUF_X1 U17 ( .A(n24), .Z(n184) );
  BUF_X2 U18 ( .A(n22), .Z(n192) );
  CLKBUF_X1 U19 ( .A(n68), .Z(n90) );
  CLKBUF_X1 U20 ( .A(n63), .Z(n76) );
  BUF_X1 U21 ( .A(n62), .Z(n81) );
  INV_X1 U22 ( .A(n65), .ZN(n64) );
  AND2_X1 U23 ( .A1(a[4]), .A2(b[4]), .ZN(shiftedA_4__8_) );
  CLKBUF_X1 U24 ( .A(n83), .Z(n65) );
  AND2_X1 U25 ( .A1(a[2]), .A2(b[6]), .ZN(shiftedA_6__8_) );
  BUF_X2 U26 ( .A(n73), .Z(n181) );
  CLKBUF_X1 U27 ( .A(a[4]), .Z(n66) );
  INV_X1 U28 ( .A(b[0]), .ZN(n67) );
  INV_X1 U29 ( .A(b[0]), .ZN(n62) );
  INV_X1 U30 ( .A(b[4]), .ZN(n68) );
  AND2_X1 U31 ( .A1(a[5]), .A2(b[1]), .ZN(shiftedA_1__6_) );
  AND2_X1 U32 ( .A1(a[2]), .A2(b[4]), .ZN(shiftedA_4__6_) );
  INV_X1 U33 ( .A(b[4]), .ZN(n58) );
  INV_X1 U34 ( .A(n88), .ZN(n69) );
  BUF_X2 U35 ( .A(n59), .Z(n88) );
  BUF_X2 U36 ( .A(n27), .Z(n180) );
  INV_X1 U37 ( .A(n89), .ZN(n70) );
  CLKBUF_X1 U38 ( .A(b[0]), .Z(n71) );
  AND2_X1 U39 ( .A1(a[6]), .A2(b[1]), .ZN(shiftedA_1__7_) );
  INV_X1 U40 ( .A(b[1]), .ZN(n61) );
  INV_X1 U41 ( .A(a[2]), .ZN(n72) );
  BUF_X2 U42 ( .A(n23), .Z(n188) );
  CLKBUF_X1 U43 ( .A(n49), .Z(n116) );
  CLKBUF_X1 U44 ( .A(n51), .Z(n109) );
  CLKBUF_X1 U45 ( .A(n50), .Z(n112) );
  CLKBUF_X1 U46 ( .A(n49), .Z(n115) );
  CLKBUF_X1 U47 ( .A(n53), .Z(n104) );
  BUF_X2 U48 ( .A(n53), .Z(n103) );
  CLKBUF_X1 U49 ( .A(n22), .Z(n190) );
  CLKBUF_X1 U50 ( .A(n18), .Z(n202) );
  CLKBUF_X1 U51 ( .A(n21), .Z(n193) );
  CLKBUF_X1 U52 ( .A(n17), .Z(n205) );
  CLKBUF_X1 U53 ( .A(n20), .Z(n196) );
  CLKBUF_X1 U54 ( .A(n19), .Z(n199) );
  BUF_X2 U55 ( .A(n57), .Z(n91) );
  BUF_X2 U56 ( .A(n60), .Z(n84) );
  BUF_X2 U57 ( .A(n56), .Z(n94) );
  BUF_X2 U58 ( .A(n55), .Z(n97) );
  CLKBUF_X1 U59 ( .A(n57), .Z(n92) );
  CLKBUF_X1 U60 ( .A(n60), .Z(n85) );
  CLKBUF_X1 U61 ( .A(n56), .Z(n95) );
  CLKBUF_X1 U62 ( .A(n55), .Z(n98) );
  CLKBUF_X1 U63 ( .A(n50), .Z(n113) );
  CLKBUF_X1 U64 ( .A(n54), .Z(n101) );
  CLKBUF_X1 U65 ( .A(n51), .Z(n110) );
  CLKBUF_X1 U66 ( .A(n52), .Z(n107) );
  CLKBUF_X1 U67 ( .A(n30), .Z(n174) );
  CLKBUF_X1 U68 ( .A(n63), .Z(n176) );
  CLKBUF_X1 U69 ( .A(n28), .Z(n178) );
  CLKBUF_X1 U70 ( .A(n56), .Z(n96) );
  CLKBUF_X1 U71 ( .A(n55), .Z(n99) );
  CLKBUF_X1 U72 ( .A(n60), .Z(n86) );
  CLKBUF_X1 U73 ( .A(n57), .Z(n93) );
  CLKBUF_X1 U74 ( .A(n54), .Z(n102) );
  CLKBUF_X1 U75 ( .A(n31), .Z(n170) );
  BUF_X1 U76 ( .A(n23), .Z(n187) );
  BUF_X1 U77 ( .A(n24), .Z(n185) );
  BUF_X1 U78 ( .A(shiftedA_54__63_), .Z(n317) );
  BUF_X1 U79 ( .A(shiftedA_53__63_), .Z(n315) );
  CLKBUF_X1 U80 ( .A(n52), .Z(n106) );
  BUF_X1 U81 ( .A(shiftedA_9__63_), .Z(n261) );
  BUF_X1 U82 ( .A(shiftedA_10__63_), .Z(n263) );
  BUF_X1 U83 ( .A(shiftedA_52__63_), .Z(n313) );
  BUF_X1 U84 ( .A(shiftedA_11__63_), .Z(n265) );
  AND2_X1 U85 ( .A1(n371), .A2(a[21]), .ZN(shiftedA_42__63_) );
  AND2_X1 U86 ( .A1(b[21]), .A2(n374), .ZN(shiftedA_21__63_) );
  AND2_X1 U87 ( .A1(n371), .A2(a[22]), .ZN(shiftedA_41__63_) );
  AND2_X1 U88 ( .A1(n371), .A2(a[23]), .ZN(shiftedA_40__63_) );
  AND2_X1 U89 ( .A1(b[23]), .A2(n374), .ZN(shiftedA_23__63_) );
  INV_X1 U90 ( .A(a[5]), .ZN(n73) );
  NOR2_X1 U91 ( .A1(n182), .A2(n129), .ZN(shiftedA_17__23_) );
  NOR2_X1 U92 ( .A1(n182), .A2(n138), .ZN(shiftedA_20__26_) );
  NOR2_X1 U93 ( .A1(n182), .A2(n147), .ZN(shiftedA_23__29_) );
  NOR2_X1 U94 ( .A1(n182), .A2(n132), .ZN(shiftedA_18__24_) );
  NOR2_X1 U95 ( .A1(n182), .A2(n141), .ZN(shiftedA_21__27_) );
  NOR2_X1 U96 ( .A1(n182), .A2(n126), .ZN(shiftedA_16__22_) );
  NOR2_X1 U97 ( .A1(n182), .A2(n135), .ZN(shiftedA_19__25_) );
  NOR2_X1 U98 ( .A1(n182), .A2(n144), .ZN(shiftedA_22__28_) );
  NOR2_X1 U99 ( .A1(n214), .A2(n89), .ZN(shiftedA_4__21_) );
  NOR2_X1 U100 ( .A1(n211), .A2(n89), .ZN(shiftedA_4__20_) );
  NOR2_X1 U101 ( .A1(n217), .A2(n89), .ZN(shiftedA_4__22_) );
  NOR2_X1 U102 ( .A1(n208), .A2(n89), .ZN(shiftedA_4__19_) );
  NOR2_X1 U103 ( .A1(n202), .A2(n89), .ZN(shiftedA_4__17_) );
  NOR2_X1 U104 ( .A1(n205), .A2(n89), .ZN(shiftedA_4__18_) );
  NOR2_X1 U105 ( .A1(n220), .A2(n89), .ZN(shiftedA_4__23_) );
  NOR2_X1 U106 ( .A1(n223), .A2(n89), .ZN(shiftedA_4__24_) );
  NOR2_X1 U107 ( .A1(n226), .A2(n89), .ZN(shiftedA_4__25_) );
  NOR2_X1 U108 ( .A1(n229), .A2(n89), .ZN(shiftedA_4__26_) );
  NOR2_X1 U109 ( .A1(n232), .A2(n89), .ZN(shiftedA_4__27_) );
  NOR2_X1 U110 ( .A1(n235), .A2(n89), .ZN(shiftedA_4__28_) );
  NOR2_X1 U111 ( .A1(n180), .A2(n138), .ZN(shiftedA_20__24_) );
  NOR2_X1 U112 ( .A1(n180), .A2(n117), .ZN(shiftedA_13__17_) );
  NOR2_X1 U113 ( .A1(n180), .A2(n126), .ZN(shiftedA_16__20_) );
  BUF_X1 U114 ( .A(n172), .Z(n173) );
  NOR2_X1 U115 ( .A1(n105), .A2(n180), .ZN(shiftedA_9__13_) );
  NOR2_X1 U116 ( .A1(n78), .A2(n120), .ZN(shiftedA_14__20_) );
  NOR2_X1 U117 ( .A1(n78), .A2(n123), .ZN(shiftedA_15__21_) );
  NOR2_X1 U118 ( .A1(n78), .A2(n117), .ZN(shiftedA_13__19_) );
  NOR2_X1 U119 ( .A1(n171), .A2(n111), .ZN(shiftedA_11__11_) );
  NOR2_X1 U120 ( .A1(n174), .A2(n111), .ZN(shiftedA_11__12_) );
  NOR2_X1 U121 ( .A1(n171), .A2(n120), .ZN(shiftedA_14__14_) );
  NOR2_X1 U122 ( .A1(n174), .A2(n120), .ZN(shiftedA_14__15_) );
  NOR2_X1 U123 ( .A1(n195), .A2(n110), .ZN(shiftedA_11__21_) );
  NOR2_X1 U124 ( .A1(n198), .A2(n110), .ZN(shiftedA_11__22_) );
  NOR2_X1 U125 ( .A1(n201), .A2(n110), .ZN(shiftedA_11__23_) );
  NOR2_X1 U126 ( .A1(n204), .A2(n110), .ZN(shiftedA_11__24_) );
  NOR2_X1 U127 ( .A1(n195), .A2(n119), .ZN(shiftedA_14__24_) );
  NOR2_X1 U128 ( .A1(n207), .A2(n110), .ZN(shiftedA_11__25_) );
  NOR2_X1 U129 ( .A1(n198), .A2(n119), .ZN(shiftedA_14__25_) );
  NOR2_X1 U130 ( .A1(n210), .A2(n110), .ZN(shiftedA_11__26_) );
  NOR2_X1 U131 ( .A1(n201), .A2(n119), .ZN(shiftedA_14__26_) );
  NOR2_X1 U132 ( .A1(n213), .A2(n110), .ZN(shiftedA_11__27_) );
  NOR2_X1 U133 ( .A1(n204), .A2(n119), .ZN(shiftedA_14__27_) );
  NOR2_X1 U134 ( .A1(n216), .A2(n110), .ZN(shiftedA_11__28_) );
  NOR2_X1 U135 ( .A1(n207), .A2(n119), .ZN(shiftedA_14__28_) );
  NOR2_X1 U136 ( .A1(n178), .A2(n141), .ZN(shiftedA_21__24_) );
  NOR2_X1 U137 ( .A1(n171), .A2(n114), .ZN(shiftedA_12__12_) );
  NOR2_X1 U138 ( .A1(n225), .A2(n80), .ZN(shiftedA_0__20_) );
  NOR2_X1 U139 ( .A1(n213), .A2(n80), .ZN(shiftedA_0__16_) );
  NOR2_X1 U140 ( .A1(n195), .A2(n81), .ZN(shiftedA_0__10_) );
  NOR2_X1 U141 ( .A1(n219), .A2(n80), .ZN(shiftedA_0__18_) );
  NOR2_X1 U142 ( .A1(n198), .A2(n81), .ZN(shiftedA_0__11_) );
  NOR2_X1 U143 ( .A1(n222), .A2(n80), .ZN(shiftedA_0__19_) );
  NOR2_X1 U144 ( .A1(n174), .A2(n114), .ZN(shiftedA_12__13_) );
  NOR2_X1 U145 ( .A1(n174), .A2(n80), .ZN(shiftedA_0__1_) );
  NOR2_X1 U146 ( .A1(n201), .A2(n81), .ZN(shiftedA_0__12_) );
  NOR2_X1 U147 ( .A1(n204), .A2(n81), .ZN(shiftedA_0__13_) );
  NOR2_X1 U148 ( .A1(n216), .A2(n80), .ZN(shiftedA_0__17_) );
  NOR2_X1 U149 ( .A1(n207), .A2(n81), .ZN(shiftedA_0__14_) );
  NOR2_X1 U150 ( .A1(n171), .A2(n123), .ZN(shiftedA_15__15_) );
  NOR2_X1 U151 ( .A1(n210), .A2(n81), .ZN(shiftedA_0__15_) );
  NOR2_X1 U152 ( .A1(n174), .A2(n123), .ZN(shiftedA_15__16_) );
  NOR2_X1 U153 ( .A1(n228), .A2(n80), .ZN(shiftedA_0__21_) );
  NOR2_X1 U154 ( .A1(n231), .A2(n80), .ZN(shiftedA_0__22_) );
  NOR2_X1 U155 ( .A1(n195), .A2(n113), .ZN(shiftedA_12__22_) );
  NOR2_X1 U156 ( .A1(n234), .A2(n80), .ZN(shiftedA_0__23_) );
  NOR2_X1 U157 ( .A1(n198), .A2(n113), .ZN(shiftedA_12__23_) );
  NOR2_X1 U158 ( .A1(n237), .A2(n80), .ZN(shiftedA_0__24_) );
  NOR2_X1 U159 ( .A1(n201), .A2(n113), .ZN(shiftedA_12__24_) );
  NOR2_X1 U160 ( .A1(n240), .A2(n80), .ZN(shiftedA_0__25_) );
  NOR2_X1 U161 ( .A1(n204), .A2(n113), .ZN(shiftedA_12__25_) );
  NOR2_X1 U162 ( .A1(n195), .A2(n122), .ZN(shiftedA_15__25_) );
  NOR2_X1 U163 ( .A1(n243), .A2(n80), .ZN(shiftedA_0__26_) );
  NOR2_X1 U164 ( .A1(n207), .A2(n113), .ZN(shiftedA_12__26_) );
  NOR2_X1 U165 ( .A1(n198), .A2(n122), .ZN(shiftedA_15__26_) );
  NOR2_X1 U166 ( .A1(n210), .A2(n113), .ZN(shiftedA_12__27_) );
  NOR2_X1 U167 ( .A1(n201), .A2(n122), .ZN(shiftedA_15__27_) );
  NOR2_X1 U168 ( .A1(n213), .A2(n113), .ZN(shiftedA_12__28_) );
  NOR2_X1 U169 ( .A1(n204), .A2(n122), .ZN(shiftedA_15__28_) );
  NOR2_X1 U170 ( .A1(n216), .A2(n113), .ZN(shiftedA_12__29_) );
  NOR2_X1 U171 ( .A1(n219), .A2(n113), .ZN(shiftedA_12__30_) );
  NOR2_X1 U172 ( .A1(n184), .A2(n93), .ZN(shiftedA_5__12_) );
  NOR2_X1 U173 ( .A1(n184), .A2(n96), .ZN(shiftedA_6__13_) );
  NOR2_X1 U174 ( .A1(n184), .A2(n131), .ZN(shiftedA_18__25_) );
  NOR2_X1 U175 ( .A1(n77), .A2(n137), .ZN(shiftedA_20__27_) );
  NOR2_X1 U176 ( .A1(n192), .A2(n110), .ZN(shiftedA_11__20_) );
  NOR2_X1 U177 ( .A1(n192), .A2(n119), .ZN(shiftedA_14__23_) );
  NOR2_X1 U178 ( .A1(n192), .A2(n113), .ZN(shiftedA_12__21_) );
  NOR2_X1 U179 ( .A1(n192), .A2(n122), .ZN(shiftedA_15__24_) );
  NOR2_X1 U180 ( .A1(n178), .A2(n117), .ZN(shiftedA_13__16_) );
  NOR2_X1 U181 ( .A1(n178), .A2(n126), .ZN(shiftedA_16__19_) );
  NOR2_X1 U182 ( .A1(n185), .A2(n88), .ZN(shiftedA_3__10_) );
  NOR2_X1 U183 ( .A1(n188), .A2(n88), .ZN(shiftedA_3__11_) );
  NOR2_X1 U184 ( .A1(n190), .A2(n87), .ZN(shiftedA_3__12_) );
  NOR2_X1 U185 ( .A1(n196), .A2(n87), .ZN(shiftedA_3__14_) );
  NOR2_X1 U186 ( .A1(n214), .A2(n87), .ZN(shiftedA_3__20_) );
  NOR2_X1 U187 ( .A1(n220), .A2(n87), .ZN(shiftedA_3__22_) );
  NOR2_X1 U188 ( .A1(n229), .A2(n88), .ZN(shiftedA_3__25_) );
  NOR2_X1 U189 ( .A1(n238), .A2(n87), .ZN(shiftedA_3__28_) );
  NOR2_X1 U190 ( .A1(n174), .A2(n108), .ZN(shiftedA_10__11_) );
  NOR2_X1 U191 ( .A1(n171), .A2(n117), .ZN(shiftedA_13__13_) );
  NOR2_X1 U192 ( .A1(n174), .A2(n117), .ZN(shiftedA_13__14_) );
  NOR2_X1 U193 ( .A1(n195), .A2(n107), .ZN(shiftedA_10__20_) );
  NOR2_X1 U194 ( .A1(n198), .A2(n107), .ZN(shiftedA_10__21_) );
  NOR2_X1 U195 ( .A1(n201), .A2(n107), .ZN(shiftedA_10__22_) );
  NOR2_X1 U196 ( .A1(n204), .A2(n107), .ZN(shiftedA_10__23_) );
  NOR2_X1 U197 ( .A1(n195), .A2(n116), .ZN(shiftedA_13__23_) );
  NOR2_X1 U198 ( .A1(n207), .A2(n107), .ZN(shiftedA_10__24_) );
  NOR2_X1 U199 ( .A1(n198), .A2(n116), .ZN(shiftedA_13__24_) );
  NOR2_X1 U200 ( .A1(n210), .A2(n107), .ZN(shiftedA_10__25_) );
  NOR2_X1 U201 ( .A1(n201), .A2(n116), .ZN(shiftedA_13__25_) );
  NOR2_X1 U202 ( .A1(n213), .A2(n107), .ZN(shiftedA_10__26_) );
  NOR2_X1 U203 ( .A1(n204), .A2(n116), .ZN(shiftedA_13__26_) );
  NOR2_X1 U204 ( .A1(n216), .A2(n107), .ZN(shiftedA_10__27_) );
  NOR2_X1 U205 ( .A1(n207), .A2(n116), .ZN(shiftedA_13__27_) );
  NOR2_X1 U206 ( .A1(n219), .A2(n107), .ZN(shiftedA_10__28_) );
  NOR2_X1 U207 ( .A1(n210), .A2(n116), .ZN(shiftedA_13__28_) );
  NOR2_X1 U208 ( .A1(n222), .A2(n106), .ZN(shiftedA_10__29_) );
  NOR2_X1 U209 ( .A1(n213), .A2(n116), .ZN(shiftedA_13__29_) );
  NOR2_X1 U210 ( .A1(n225), .A2(n106), .ZN(shiftedA_10__30_) );
  NOR2_X1 U211 ( .A1(n216), .A2(n116), .ZN(shiftedA_13__30_) );
  NOR2_X1 U212 ( .A1(n184), .A2(n99), .ZN(shiftedA_7__14_) );
  NOR2_X1 U213 ( .A1(n184), .A2(n134), .ZN(shiftedA_19__26_) );
  NOR2_X1 U214 ( .A1(n76), .A2(n120), .ZN(shiftedA_14__16_) );
  NOR2_X1 U215 ( .A1(n76), .A2(n129), .ZN(shiftedA_17__19_) );
  NOR2_X1 U216 ( .A1(n76), .A2(n138), .ZN(shiftedA_20__22_) );
  NOR2_X1 U217 ( .A1(n76), .A2(n147), .ZN(shiftedA_23__25_) );
  NOR2_X1 U218 ( .A1(n77), .A2(n125), .ZN(shiftedA_16__23_) );
  NOR2_X1 U219 ( .A1(n192), .A2(n107), .ZN(shiftedA_10__19_) );
  NOR2_X1 U220 ( .A1(n192), .A2(n116), .ZN(shiftedA_13__22_) );
  NOR2_X1 U221 ( .A1(n63), .A2(n108), .ZN(shiftedA_10__12_) );
  NOR2_X1 U222 ( .A1(n105), .A2(n178), .ZN(shiftedA_9__12_) );
  NOR2_X1 U223 ( .A1(n105), .A2(n77), .ZN(shiftedA_9__16_) );
  NOR2_X1 U224 ( .A1(n105), .A2(n78), .ZN(shiftedA_9__15_) );
  NOR2_X1 U225 ( .A1(n76), .A2(n132), .ZN(shiftedA_18__20_) );
  NOR2_X1 U226 ( .A1(n76), .A2(n141), .ZN(shiftedA_21__23_) );
  NOR2_X1 U227 ( .A1(n76), .A2(n150), .ZN(shiftedA_24__26_) );
  NOR2_X1 U228 ( .A1(n190), .A2(n86), .ZN(shiftedA_2__11_) );
  NOR2_X1 U229 ( .A1(n193), .A2(n86), .ZN(shiftedA_2__12_) );
  NOR2_X1 U230 ( .A1(n196), .A2(n86), .ZN(shiftedA_2__13_) );
  NOR2_X1 U231 ( .A1(n199), .A2(n86), .ZN(shiftedA_2__14_) );
  NOR2_X1 U232 ( .A1(n202), .A2(n86), .ZN(shiftedA_2__15_) );
  NOR2_X1 U233 ( .A1(n205), .A2(n86), .ZN(shiftedA_2__16_) );
  NOR2_X1 U234 ( .A1(n78), .A2(n93), .ZN(shiftedA_5__11_) );
  NOR2_X1 U235 ( .A1(n170), .A2(n129), .ZN(shiftedA_17__17_) );
  NOR2_X1 U236 ( .A1(n173), .A2(n129), .ZN(shiftedA_17__18_) );
  NOR2_X1 U237 ( .A1(n63), .A2(n111), .ZN(shiftedA_11__13_) );
  NOR2_X1 U238 ( .A1(n183), .A2(n111), .ZN(shiftedA_11__17_) );
  NOR2_X1 U239 ( .A1(n187), .A2(n93), .ZN(shiftedA_5__13_) );
  NOR2_X1 U240 ( .A1(n177), .A2(n111), .ZN(shiftedA_11__14_) );
  NOR2_X1 U241 ( .A1(n190), .A2(n93), .ZN(shiftedA_5__14_) );
  NOR2_X1 U242 ( .A1(n179), .A2(n111), .ZN(shiftedA_11__15_) );
  NOR2_X1 U243 ( .A1(n193), .A2(n93), .ZN(shiftedA_5__15_) );
  NOR2_X1 U244 ( .A1(n196), .A2(n93), .ZN(shiftedA_5__16_) );
  NOR2_X1 U245 ( .A1(n177), .A2(n129), .ZN(shiftedA_17__20_) );
  NOR2_X1 U246 ( .A1(n170), .A2(n138), .ZN(shiftedA_20__20_) );
  NOR2_X1 U247 ( .A1(n179), .A2(n129), .ZN(shiftedA_17__21_) );
  NOR2_X1 U248 ( .A1(n173), .A2(n138), .ZN(shiftedA_20__21_) );
  NOR2_X1 U249 ( .A1(n170), .A2(n147), .ZN(shiftedA_23__23_) );
  NOR2_X1 U250 ( .A1(n177), .A2(n138), .ZN(shiftedA_20__23_) );
  NOR2_X1 U251 ( .A1(n173), .A2(n147), .ZN(shiftedA_23__24_) );
  NOR2_X1 U252 ( .A1(n177), .A2(n147), .ZN(shiftedA_23__26_) );
  NOR2_X1 U253 ( .A1(n170), .A2(n156), .ZN(shiftedA_26__26_) );
  NOR2_X1 U254 ( .A1(n179), .A2(n147), .ZN(shiftedA_23__27_) );
  NOR2_X1 U255 ( .A1(n173), .A2(n156), .ZN(shiftedA_26__27_) );
  NOR2_X1 U256 ( .A1(n190), .A2(n96), .ZN(shiftedA_6__15_) );
  NOR2_X1 U257 ( .A1(n179), .A2(n96), .ZN(shiftedA_6__10_) );
  NOR2_X1 U258 ( .A1(n26), .A2(n123), .ZN(shiftedA_15__17_) );
  NOR2_X1 U259 ( .A1(n182), .A2(n96), .ZN(shiftedA_6__12_) );
  NOR2_X1 U260 ( .A1(n177), .A2(n123), .ZN(shiftedA_15__18_) );
  NOR2_X1 U261 ( .A1(n188), .A2(n96), .ZN(shiftedA_6__14_) );
  NOR2_X1 U262 ( .A1(n193), .A2(n96), .ZN(shiftedA_6__16_) );
  NOR2_X1 U263 ( .A1(n179), .A2(n123), .ZN(shiftedA_15__19_) );
  NOR2_X1 U264 ( .A1(n170), .A2(n141), .ZN(shiftedA_21__21_) );
  NOR2_X1 U265 ( .A1(n173), .A2(n141), .ZN(shiftedA_21__22_) );
  NOR2_X1 U266 ( .A1(n179), .A2(n141), .ZN(shiftedA_21__25_) );
  NOR2_X1 U267 ( .A1(n187), .A2(n102), .ZN(shiftedA_8__16_) );
  NOR2_X1 U268 ( .A1(n177), .A2(n102), .ZN(shiftedA_8__11_) );
  NOR2_X1 U269 ( .A1(n179), .A2(n102), .ZN(shiftedA_8__12_) );
  NOR2_X1 U270 ( .A1(n182), .A2(n102), .ZN(shiftedA_8__14_) );
  NOR2_X1 U271 ( .A1(n185), .A2(n102), .ZN(shiftedA_8__15_) );
  NOR2_X1 U272 ( .A1(n76), .A2(n117), .ZN(shiftedA_13__15_) );
  NOR2_X1 U273 ( .A1(n170), .A2(n132), .ZN(shiftedA_18__18_) );
  NOR2_X1 U274 ( .A1(n173), .A2(n132), .ZN(shiftedA_18__19_) );
  NOR2_X1 U275 ( .A1(n183), .A2(n114), .ZN(shiftedA_12__18_) );
  NOR2_X1 U276 ( .A1(n63), .A2(n114), .ZN(shiftedA_12__14_) );
  NOR2_X1 U277 ( .A1(n170), .A2(n150), .ZN(shiftedA_24__24_) );
  NOR2_X1 U278 ( .A1(n173), .A2(n150), .ZN(shiftedA_24__25_) );
  NOR2_X1 U279 ( .A1(n169), .A2(n159), .ZN(shiftedA_27__27_) );
  NOR2_X1 U280 ( .A1(n169), .A2(n168), .ZN(shiftedA_30__30_) );
  NOR2_X1 U281 ( .A1(n191), .A2(n83), .ZN(shiftedA_1__10_) );
  NOR2_X1 U282 ( .A1(n199), .A2(n68), .ZN(shiftedA_4__16_) );
  NOR2_X1 U283 ( .A1(n209), .A2(n65), .ZN(shiftedA_1__16_) );
  NOR2_X1 U284 ( .A1(n183), .A2(n68), .ZN(shiftedA_4__10_) );
  NOR2_X1 U285 ( .A1(n194), .A2(n83), .ZN(shiftedA_1__11_) );
  NOR2_X1 U286 ( .A1(n185), .A2(n68), .ZN(shiftedA_4__11_) );
  NOR2_X1 U287 ( .A1(n197), .A2(n83), .ZN(shiftedA_1__12_) );
  NOR2_X1 U288 ( .A1(n187), .A2(n68), .ZN(shiftedA_4__12_) );
  NOR2_X1 U289 ( .A1(n200), .A2(n83), .ZN(shiftedA_1__13_) );
  NOR2_X1 U290 ( .A1(n190), .A2(n68), .ZN(shiftedA_4__13_) );
  NOR2_X1 U291 ( .A1(n203), .A2(n83), .ZN(shiftedA_1__14_) );
  NOR2_X1 U292 ( .A1(n193), .A2(n68), .ZN(shiftedA_4__14_) );
  NOR2_X1 U293 ( .A1(n206), .A2(n65), .ZN(shiftedA_1__15_) );
  NOR2_X1 U294 ( .A1(n196), .A2(n68), .ZN(shiftedA_4__15_) );
  NOR2_X1 U295 ( .A1(n187), .A2(n99), .ZN(shiftedA_7__15_) );
  NOR2_X1 U296 ( .A1(n177), .A2(n99), .ZN(shiftedA_7__10_) );
  NOR2_X1 U297 ( .A1(n179), .A2(n99), .ZN(shiftedA_7__11_) );
  NOR2_X1 U298 ( .A1(n173), .A2(n126), .ZN(shiftedA_16__17_) );
  NOR2_X1 U299 ( .A1(n26), .A2(n126), .ZN(shiftedA_16__18_) );
  NOR2_X1 U300 ( .A1(n182), .A2(n99), .ZN(shiftedA_7__13_) );
  NOR2_X1 U301 ( .A1(n170), .A2(n126), .ZN(shiftedA_16__16_) );
  NOR2_X1 U302 ( .A1(n190), .A2(n99), .ZN(shiftedA_7__16_) );
  NOR2_X1 U303 ( .A1(n170), .A2(n153), .ZN(shiftedA_25__25_) );
  NOR2_X1 U304 ( .A1(n173), .A2(n153), .ZN(shiftedA_25__26_) );
  NOR2_X1 U305 ( .A1(n26), .A2(n153), .ZN(shiftedA_25__27_) );
  NOR2_X1 U306 ( .A1(n179), .A2(n91), .ZN(shiftedA_5__9_) );
  NOR2_X1 U307 ( .A1(n208), .A2(n85), .ZN(shiftedA_2__17_) );
  NOR2_X1 U308 ( .A1(n202), .A2(n92), .ZN(shiftedA_5__18_) );
  NOR2_X1 U309 ( .A1(n211), .A2(n85), .ZN(shiftedA_2__18_) );
  NOR2_X1 U310 ( .A1(n190), .A2(n101), .ZN(shiftedA_8__17_) );
  NOR2_X1 U311 ( .A1(n199), .A2(n92), .ZN(shiftedA_5__17_) );
  NOR2_X1 U312 ( .A1(n193), .A2(n101), .ZN(shiftedA_8__18_) );
  NOR2_X1 U313 ( .A1(n205), .A2(n92), .ZN(shiftedA_5__19_) );
  NOR2_X1 U314 ( .A1(n214), .A2(n85), .ZN(shiftedA_2__19_) );
  NOR2_X1 U315 ( .A1(n196), .A2(n101), .ZN(shiftedA_8__19_) );
  NOR2_X1 U316 ( .A1(n208), .A2(n92), .ZN(shiftedA_5__20_) );
  NOR2_X1 U317 ( .A1(n217), .A2(n85), .ZN(shiftedA_2__20_) );
  NOR2_X1 U318 ( .A1(n199), .A2(n101), .ZN(shiftedA_8__20_) );
  NOR2_X1 U319 ( .A1(n211), .A2(n92), .ZN(shiftedA_5__21_) );
  NOR2_X1 U320 ( .A1(n220), .A2(n85), .ZN(shiftedA_2__21_) );
  NOR2_X1 U321 ( .A1(n202), .A2(n101), .ZN(shiftedA_8__21_) );
  NOR2_X1 U322 ( .A1(n214), .A2(n92), .ZN(shiftedA_5__22_) );
  NOR2_X1 U323 ( .A1(n223), .A2(n85), .ZN(shiftedA_2__22_) );
  NOR2_X1 U324 ( .A1(n205), .A2(n101), .ZN(shiftedA_8__22_) );
  NOR2_X1 U325 ( .A1(n217), .A2(n92), .ZN(shiftedA_5__23_) );
  NOR2_X1 U326 ( .A1(n226), .A2(n85), .ZN(shiftedA_2__23_) );
  NOR2_X1 U327 ( .A1(n208), .A2(n101), .ZN(shiftedA_8__23_) );
  NOR2_X1 U328 ( .A1(n220), .A2(n92), .ZN(shiftedA_5__24_) );
  NOR2_X1 U329 ( .A1(n229), .A2(n85), .ZN(shiftedA_2__24_) );
  NOR2_X1 U330 ( .A1(n211), .A2(n101), .ZN(shiftedA_8__24_) );
  NOR2_X1 U331 ( .A1(n223), .A2(n92), .ZN(shiftedA_5__25_) );
  NOR2_X1 U332 ( .A1(n232), .A2(n85), .ZN(shiftedA_2__25_) );
  NOR2_X1 U333 ( .A1(n214), .A2(n101), .ZN(shiftedA_8__25_) );
  NOR2_X1 U334 ( .A1(n226), .A2(n92), .ZN(shiftedA_5__26_) );
  NOR2_X1 U335 ( .A1(n235), .A2(n85), .ZN(shiftedA_2__26_) );
  NOR2_X1 U336 ( .A1(n217), .A2(n101), .ZN(shiftedA_8__26_) );
  NOR2_X1 U337 ( .A1(n191), .A2(n128), .ZN(shiftedA_17__26_) );
  NOR2_X1 U338 ( .A1(n229), .A2(n92), .ZN(shiftedA_5__27_) );
  NOR2_X1 U339 ( .A1(n220), .A2(n101), .ZN(shiftedA_8__27_) );
  NOR2_X1 U340 ( .A1(n194), .A2(n128), .ZN(shiftedA_17__27_) );
  NOR2_X1 U341 ( .A1(n232), .A2(n92), .ZN(shiftedA_5__28_) );
  NOR2_X1 U342 ( .A1(n188), .A2(n128), .ZN(shiftedA_17__25_) );
  NOR2_X1 U343 ( .A1(n238), .A2(n85), .ZN(shiftedA_2__27_) );
  NOR2_X1 U344 ( .A1(n169), .A2(n84), .ZN(shiftedA_2__2_) );
  NOR2_X1 U345 ( .A1(n169), .A2(n100), .ZN(shiftedA_8__8_) );
  NOR2_X1 U346 ( .A1(n241), .A2(n85), .ZN(shiftedA_2__28_) );
  NOR2_X1 U347 ( .A1(n244), .A2(n84), .ZN(shiftedA_2__29_) );
  NOR2_X1 U348 ( .A1(n185), .A2(n84), .ZN(shiftedA_2__9_) );
  NOR2_X1 U349 ( .A1(n185), .A2(n128), .ZN(shiftedA_17__24_) );
  NOR2_X1 U350 ( .A1(n211), .A2(n88), .ZN(shiftedA_3__19_) );
  NOR2_X1 U351 ( .A1(n208), .A2(n87), .ZN(shiftedA_3__18_) );
  NOR2_X1 U352 ( .A1(n202), .A2(n87), .ZN(shiftedA_3__16_) );
  NOR2_X1 U353 ( .A1(n104), .A2(n193), .ZN(shiftedA_9__19_) );
  NOR2_X1 U354 ( .A1(n199), .A2(n95), .ZN(shiftedA_6__18_) );
  NOR2_X1 U355 ( .A1(n193), .A2(n88), .ZN(shiftedA_3__13_) );
  NOR2_X1 U356 ( .A1(n196), .A2(n95), .ZN(shiftedA_6__17_) );
  NOR2_X1 U357 ( .A1(n104), .A2(n190), .ZN(shiftedA_9__18_) );
  NOR2_X1 U358 ( .A1(n199), .A2(n88), .ZN(shiftedA_3__15_) );
  NOR2_X1 U359 ( .A1(n205), .A2(n88), .ZN(shiftedA_3__17_) );
  NOR2_X1 U360 ( .A1(n104), .A2(n188), .ZN(shiftedA_9__17_) );
  NOR2_X1 U361 ( .A1(n202), .A2(n95), .ZN(shiftedA_6__19_) );
  NOR2_X1 U362 ( .A1(n104), .A2(n196), .ZN(shiftedA_9__20_) );
  NOR2_X1 U363 ( .A1(n205), .A2(n95), .ZN(shiftedA_6__20_) );
  NOR2_X1 U364 ( .A1(n217), .A2(n88), .ZN(shiftedA_3__21_) );
  NOR2_X1 U365 ( .A1(n104), .A2(n199), .ZN(shiftedA_9__21_) );
  NOR2_X1 U366 ( .A1(n208), .A2(n95), .ZN(shiftedA_6__21_) );
  NOR2_X1 U367 ( .A1(n104), .A2(n202), .ZN(shiftedA_9__22_) );
  NOR2_X1 U368 ( .A1(n211), .A2(n95), .ZN(shiftedA_6__22_) );
  NOR2_X1 U369 ( .A1(n223), .A2(n88), .ZN(shiftedA_3__23_) );
  NOR2_X1 U370 ( .A1(n104), .A2(n205), .ZN(shiftedA_9__23_) );
  NOR2_X1 U371 ( .A1(n214), .A2(n95), .ZN(shiftedA_6__23_) );
  NOR2_X1 U372 ( .A1(n226), .A2(n87), .ZN(shiftedA_3__24_) );
  NOR2_X1 U373 ( .A1(n104), .A2(n208), .ZN(shiftedA_9__24_) );
  NOR2_X1 U374 ( .A1(n217), .A2(n95), .ZN(shiftedA_6__24_) );
  NOR2_X1 U375 ( .A1(n104), .A2(n211), .ZN(shiftedA_9__25_) );
  NOR2_X1 U376 ( .A1(n220), .A2(n95), .ZN(shiftedA_6__25_) );
  NOR2_X1 U377 ( .A1(n232), .A2(n87), .ZN(shiftedA_3__26_) );
  NOR2_X1 U378 ( .A1(n104), .A2(n214), .ZN(shiftedA_9__26_) );
  NOR2_X1 U379 ( .A1(n223), .A2(n95), .ZN(shiftedA_6__26_) );
  NOR2_X1 U380 ( .A1(n235), .A2(n88), .ZN(shiftedA_3__27_) );
  NOR2_X1 U381 ( .A1(n104), .A2(n217), .ZN(shiftedA_9__27_) );
  NOR2_X1 U382 ( .A1(n226), .A2(n95), .ZN(shiftedA_6__27_) );
  NOR2_X1 U383 ( .A1(n191), .A2(n131), .ZN(shiftedA_18__27_) );
  NOR2_X1 U384 ( .A1(n104), .A2(n220), .ZN(shiftedA_9__28_) );
  NOR2_X1 U385 ( .A1(n229), .A2(n95), .ZN(shiftedA_6__28_) );
  NOR2_X1 U386 ( .A1(n194), .A2(n131), .ZN(shiftedA_18__28_) );
  NOR2_X1 U387 ( .A1(n103), .A2(n223), .ZN(shiftedA_9__29_) );
  NOR2_X1 U388 ( .A1(n103), .A2(n226), .ZN(shiftedA_9__30_) );
  NOR2_X1 U389 ( .A1(n177), .A2(n94), .ZN(shiftedA_6__9_) );
  NOR2_X1 U390 ( .A1(n188), .A2(n131), .ZN(shiftedA_18__26_) );
  NOR2_X1 U391 ( .A1(n188), .A2(n140), .ZN(shiftedA_21__29_) );
  NOR2_X1 U392 ( .A1(n169), .A2(n94), .ZN(shiftedA_6__6_) );
  NOR2_X1 U393 ( .A1(n185), .A2(n140), .ZN(shiftedA_21__28_) );
  NOR2_X1 U394 ( .A1(n183), .A2(n108), .ZN(shiftedA_10__16_) );
  NOR2_X1 U395 ( .A1(n170), .A2(n135), .ZN(shiftedA_19__19_) );
  NOR2_X1 U396 ( .A1(n173), .A2(n135), .ZN(shiftedA_19__20_) );
  NOR2_X1 U397 ( .A1(n26), .A2(n135), .ZN(shiftedA_19__21_) );
  NOR2_X1 U398 ( .A1(n170), .A2(n144), .ZN(shiftedA_22__22_) );
  NOR2_X1 U399 ( .A1(n173), .A2(n144), .ZN(shiftedA_22__23_) );
  NOR2_X1 U400 ( .A1(n26), .A2(n144), .ZN(shiftedA_22__24_) );
  NOR2_X1 U401 ( .A1(n221), .A2(n82), .ZN(shiftedA_1__20_) );
  NOR2_X1 U402 ( .A1(n215), .A2(n82), .ZN(shiftedA_1__18_) );
  NOR2_X1 U403 ( .A1(n218), .A2(n82), .ZN(shiftedA_1__19_) );
  NOR2_X1 U404 ( .A1(n170), .A2(n82), .ZN(shiftedA_1__1_) );
  NOR2_X1 U405 ( .A1(n212), .A2(n82), .ZN(shiftedA_1__17_) );
  NOR2_X1 U406 ( .A1(n224), .A2(n82), .ZN(shiftedA_1__21_) );
  NOR2_X1 U407 ( .A1(n227), .A2(n82), .ZN(shiftedA_1__22_) );
  NOR2_X1 U408 ( .A1(n230), .A2(n82), .ZN(shiftedA_1__23_) );
  NOR2_X1 U409 ( .A1(n233), .A2(n82), .ZN(shiftedA_1__24_) );
  NOR2_X1 U410 ( .A1(n236), .A2(n82), .ZN(shiftedA_1__25_) );
  NOR2_X1 U411 ( .A1(n239), .A2(n82), .ZN(shiftedA_1__26_) );
  NOR2_X1 U412 ( .A1(n242), .A2(n82), .ZN(shiftedA_1__27_) );
  NOR2_X1 U413 ( .A1(n169), .A2(n162), .ZN(shiftedA_28__28_) );
  NOR2_X1 U414 ( .A1(n196), .A2(n98), .ZN(shiftedA_7__18_) );
  NOR2_X1 U415 ( .A1(n193), .A2(n98), .ZN(shiftedA_7__17_) );
  NOR2_X1 U416 ( .A1(n199), .A2(n98), .ZN(shiftedA_7__19_) );
  NOR2_X1 U417 ( .A1(n202), .A2(n98), .ZN(shiftedA_7__20_) );
  NOR2_X1 U418 ( .A1(n205), .A2(n98), .ZN(shiftedA_7__21_) );
  NOR2_X1 U419 ( .A1(n208), .A2(n98), .ZN(shiftedA_7__22_) );
  NOR2_X1 U420 ( .A1(n211), .A2(n98), .ZN(shiftedA_7__23_) );
  NOR2_X1 U421 ( .A1(n214), .A2(n98), .ZN(shiftedA_7__24_) );
  NOR2_X1 U422 ( .A1(n217), .A2(n98), .ZN(shiftedA_7__25_) );
  NOR2_X1 U423 ( .A1(n191), .A2(n125), .ZN(shiftedA_16__25_) );
  NOR2_X1 U424 ( .A1(n220), .A2(n98), .ZN(shiftedA_7__26_) );
  NOR2_X1 U425 ( .A1(n194), .A2(n125), .ZN(shiftedA_16__26_) );
  NOR2_X1 U426 ( .A1(n223), .A2(n98), .ZN(shiftedA_7__27_) );
  NOR2_X1 U427 ( .A1(n197), .A2(n125), .ZN(shiftedA_16__27_) );
  NOR2_X1 U428 ( .A1(n226), .A2(n98), .ZN(shiftedA_7__28_) );
  NOR2_X1 U429 ( .A1(n200), .A2(n125), .ZN(shiftedA_16__28_) );
  NOR2_X1 U430 ( .A1(n191), .A2(n134), .ZN(shiftedA_19__28_) );
  NOR2_X1 U431 ( .A1(n188), .A2(n125), .ZN(shiftedA_16__24_) );
  NOR2_X1 U432 ( .A1(n187), .A2(n134), .ZN(shiftedA_19__27_) );
  NOR2_X1 U433 ( .A1(n169), .A2(n97), .ZN(shiftedA_7__7_) );
  NOR2_X1 U434 ( .A1(n171), .A2(n108), .ZN(shiftedA_10__10_) );
  NOR2_X1 U435 ( .A1(n169), .A2(n103), .ZN(shiftedA_9__9_) );
  NOR2_X1 U436 ( .A1(n183), .A2(n84), .ZN(shiftedA_2__8_) );
  NOR2_X1 U437 ( .A1(n169), .A2(n91), .ZN(shiftedA_5__5_) );
  NOR2_X1 U438 ( .A1(n177), .A2(n91), .ZN(shiftedA_5__8_) );
  BUF_X2 U439 ( .A(shiftedA_58__63_), .Z(n328) );
  BUF_X2 U440 ( .A(shiftedA_56__63_), .Z(n322) );
  BUF_X2 U441 ( .A(shiftedA_58__63_), .Z(n329) );
  BUF_X2 U442 ( .A(shiftedA_56__63_), .Z(n323) );
  NOR2_X1 U443 ( .A1(n182), .A2(n156), .ZN(shiftedA_26__32_) );
  NOR2_X1 U444 ( .A1(n182), .A2(n150), .ZN(shiftedA_24__30_) );
  NOR2_X1 U445 ( .A1(n182), .A2(n153), .ZN(shiftedA_25__31_) );
  NOR2_X1 U446 ( .A1(n180), .A2(n165), .ZN(shiftedA_29__33_) );
  NOR2_X1 U447 ( .A1(n180), .A2(n159), .ZN(shiftedA_27__31_) );
  NOR2_X1 U448 ( .A1(n180), .A2(n168), .ZN(shiftedA_30__34_) );
  BUF_X1 U449 ( .A(shiftedA_58__63_), .Z(n330) );
  NOR2_X1 U450 ( .A1(n178), .A2(n165), .ZN(shiftedA_29__32_) );
  NOR2_X1 U451 ( .A1(n219), .A2(n110), .ZN(shiftedA_11__29_) );
  NOR2_X1 U452 ( .A1(n210), .A2(n119), .ZN(shiftedA_14__29_) );
  NOR2_X1 U453 ( .A1(n222), .A2(n109), .ZN(shiftedA_11__30_) );
  NOR2_X1 U454 ( .A1(n213), .A2(n119), .ZN(shiftedA_14__30_) );
  NOR2_X1 U455 ( .A1(n225), .A2(n109), .ZN(shiftedA_11__31_) );
  NOR2_X1 U456 ( .A1(n216), .A2(n119), .ZN(shiftedA_14__31_) );
  NOR2_X1 U457 ( .A1(n228), .A2(n109), .ZN(shiftedA_11__32_) );
  NOR2_X1 U458 ( .A1(n219), .A2(n119), .ZN(shiftedA_14__32_) );
  NOR2_X1 U459 ( .A1(n231), .A2(n109), .ZN(shiftedA_11__33_) );
  NOR2_X1 U460 ( .A1(n222), .A2(n118), .ZN(shiftedA_14__33_) );
  NOR2_X1 U461 ( .A1(n225), .A2(n118), .ZN(shiftedA_14__34_) );
  NOR2_X1 U462 ( .A1(n234), .A2(n109), .ZN(shiftedA_11__34_) );
  NOR2_X1 U463 ( .A1(n228), .A2(n118), .ZN(shiftedA_14__35_) );
  NOR2_X1 U464 ( .A1(n237), .A2(n109), .ZN(shiftedA_11__35_) );
  NOR2_X1 U465 ( .A1(n231), .A2(n118), .ZN(shiftedA_14__36_) );
  NOR2_X1 U466 ( .A1(n240), .A2(n109), .ZN(shiftedA_11__36_) );
  NOR2_X1 U467 ( .A1(n234), .A2(n118), .ZN(shiftedA_14__37_) );
  NOR2_X1 U468 ( .A1(n243), .A2(n109), .ZN(shiftedA_11__37_) );
  NOR2_X1 U469 ( .A1(n237), .A2(n118), .ZN(shiftedA_14__38_) );
  NOR2_X1 U470 ( .A1(n240), .A2(n118), .ZN(shiftedA_14__39_) );
  NOR2_X1 U471 ( .A1(n243), .A2(n118), .ZN(shiftedA_14__40_) );
  NOR2_X1 U472 ( .A1(n178), .A2(n159), .ZN(shiftedA_27__30_) );
  NOR2_X1 U473 ( .A1(n178), .A2(n168), .ZN(shiftedA_30__33_) );
  NOR2_X1 U474 ( .A1(n207), .A2(n122), .ZN(shiftedA_15__29_) );
  NOR2_X1 U475 ( .A1(n210), .A2(n122), .ZN(shiftedA_15__30_) );
  NOR2_X1 U476 ( .A1(n222), .A2(n112), .ZN(shiftedA_12__31_) );
  NOR2_X1 U477 ( .A1(n213), .A2(n122), .ZN(shiftedA_15__31_) );
  NOR2_X1 U478 ( .A1(n225), .A2(n112), .ZN(shiftedA_12__32_) );
  NOR2_X1 U479 ( .A1(n216), .A2(n122), .ZN(shiftedA_15__32_) );
  NOR2_X1 U480 ( .A1(n228), .A2(n112), .ZN(shiftedA_12__33_) );
  NOR2_X1 U481 ( .A1(n219), .A2(n122), .ZN(shiftedA_15__33_) );
  NOR2_X1 U482 ( .A1(n231), .A2(n112), .ZN(shiftedA_12__34_) );
  NOR2_X1 U483 ( .A1(n222), .A2(n121), .ZN(shiftedA_15__34_) );
  NOR2_X1 U484 ( .A1(n234), .A2(n112), .ZN(shiftedA_12__35_) );
  NOR2_X1 U485 ( .A1(n225), .A2(n121), .ZN(shiftedA_15__35_) );
  NOR2_X1 U486 ( .A1(n237), .A2(n112), .ZN(shiftedA_12__36_) );
  NOR2_X1 U487 ( .A1(n228), .A2(n121), .ZN(shiftedA_15__36_) );
  NOR2_X1 U488 ( .A1(n240), .A2(n112), .ZN(shiftedA_12__37_) );
  NOR2_X1 U489 ( .A1(n231), .A2(n121), .ZN(shiftedA_15__37_) );
  NOR2_X1 U490 ( .A1(n243), .A2(n112), .ZN(shiftedA_12__38_) );
  NOR2_X1 U491 ( .A1(n234), .A2(n121), .ZN(shiftedA_15__38_) );
  NOR2_X1 U492 ( .A1(n237), .A2(n121), .ZN(shiftedA_15__39_) );
  NOR2_X1 U493 ( .A1(n240), .A2(n121), .ZN(shiftedA_15__40_) );
  NOR2_X1 U494 ( .A1(n243), .A2(n121), .ZN(shiftedA_15__41_) );
  NOR2_X1 U495 ( .A1(n184), .A2(n149), .ZN(shiftedA_24__31_) );
  NOR2_X1 U496 ( .A1(n77), .A2(n164), .ZN(shiftedA_29__36_) );
  NOR2_X1 U497 ( .A1(n246), .A2(n109), .ZN(shiftedA_11__38_) );
  NOR2_X1 U498 ( .A1(n249), .A2(n109), .ZN(shiftedA_11__39_) );
  NOR2_X1 U499 ( .A1(n252), .A2(n109), .ZN(shiftedA_11__40_) );
  NOR2_X1 U500 ( .A1(n255), .A2(n109), .ZN(shiftedA_11__41_) );
  NOR2_X1 U501 ( .A1(n246), .A2(n118), .ZN(shiftedA_14__41_) );
  NOR2_X1 U502 ( .A1(n77), .A2(n167), .ZN(shiftedA_30__37_) );
  NOR2_X1 U503 ( .A1(n246), .A2(n112), .ZN(shiftedA_12__39_) );
  NOR2_X1 U504 ( .A1(n249), .A2(n112), .ZN(shiftedA_12__40_) );
  NOR2_X1 U505 ( .A1(n252), .A2(n112), .ZN(shiftedA_12__41_) );
  NOR2_X1 U506 ( .A1(n255), .A2(n112), .ZN(shiftedA_12__42_) );
  NOR2_X1 U507 ( .A1(n228), .A2(n106), .ZN(shiftedA_10__31_) );
  NOR2_X1 U508 ( .A1(n219), .A2(n116), .ZN(shiftedA_13__31_) );
  NOR2_X1 U509 ( .A1(n231), .A2(n106), .ZN(shiftedA_10__32_) );
  NOR2_X1 U510 ( .A1(n222), .A2(n115), .ZN(shiftedA_13__32_) );
  NOR2_X1 U511 ( .A1(n234), .A2(n106), .ZN(shiftedA_10__33_) );
  NOR2_X1 U512 ( .A1(n225), .A2(n115), .ZN(shiftedA_13__33_) );
  NOR2_X1 U513 ( .A1(n228), .A2(n115), .ZN(shiftedA_13__34_) );
  NOR2_X1 U514 ( .A1(n237), .A2(n106), .ZN(shiftedA_10__34_) );
  NOR2_X1 U515 ( .A1(n231), .A2(n115), .ZN(shiftedA_13__35_) );
  NOR2_X1 U516 ( .A1(n240), .A2(n106), .ZN(shiftedA_10__35_) );
  NOR2_X1 U517 ( .A1(n234), .A2(n115), .ZN(shiftedA_13__36_) );
  NOR2_X1 U518 ( .A1(n243), .A2(n106), .ZN(shiftedA_10__36_) );
  NOR2_X1 U519 ( .A1(n237), .A2(n115), .ZN(shiftedA_13__37_) );
  NOR2_X1 U520 ( .A1(n240), .A2(n115), .ZN(shiftedA_13__38_) );
  NOR2_X1 U521 ( .A1(n243), .A2(n115), .ZN(shiftedA_13__39_) );
  NOR2_X1 U522 ( .A1(n184), .A2(n143), .ZN(shiftedA_22__29_) );
  NOR2_X1 U523 ( .A1(n184), .A2(n161), .ZN(shiftedA_28__35_) );
  NOR2_X1 U524 ( .A1(n76), .A2(n156), .ZN(shiftedA_26__28_) );
  NOR2_X1 U525 ( .A1(n77), .A2(n152), .ZN(shiftedA_25__32_) );
  NOR2_X1 U526 ( .A1(n246), .A2(n106), .ZN(shiftedA_10__37_) );
  NOR2_X1 U527 ( .A1(n249), .A2(n106), .ZN(shiftedA_10__38_) );
  NOR2_X1 U528 ( .A1(n252), .A2(n106), .ZN(shiftedA_10__39_) );
  NOR2_X1 U529 ( .A1(n255), .A2(n106), .ZN(shiftedA_10__40_) );
  NOR2_X1 U530 ( .A1(n246), .A2(n115), .ZN(shiftedA_13__40_) );
  NOR2_X1 U531 ( .A1(n249), .A2(n115), .ZN(shiftedA_13__41_) );
  NOR2_X1 U532 ( .A1(n252), .A2(n115), .ZN(shiftedA_13__42_) );
  NOR2_X1 U533 ( .A1(n177), .A2(n156), .ZN(shiftedA_26__29_) );
  NOR2_X1 U534 ( .A1(n179), .A2(n156), .ZN(shiftedA_26__30_) );
  NOR2_X1 U535 ( .A1(n169), .A2(n165), .ZN(shiftedA_29__29_) );
  NOR2_X1 U536 ( .A1(n183), .A2(n165), .ZN(shiftedA_29__35_) );
  NOR2_X1 U537 ( .A1(n78), .A2(n159), .ZN(shiftedA_27__33_) );
  NOR2_X1 U538 ( .A1(n78), .A2(n168), .ZN(shiftedA_30__36_) );
  NOR2_X1 U539 ( .A1(n177), .A2(n153), .ZN(shiftedA_25__28_) );
  NOR2_X1 U540 ( .A1(n179), .A2(n153), .ZN(shiftedA_25__29_) );
  NOR2_X1 U541 ( .A1(n223), .A2(n101), .ZN(shiftedA_8__28_) );
  NOR2_X1 U542 ( .A1(n197), .A2(n128), .ZN(shiftedA_17__28_) );
  NOR2_X1 U543 ( .A1(n235), .A2(n91), .ZN(shiftedA_5__29_) );
  NOR2_X1 U544 ( .A1(n226), .A2(n100), .ZN(shiftedA_8__29_) );
  NOR2_X1 U545 ( .A1(n200), .A2(n128), .ZN(shiftedA_17__29_) );
  NOR2_X1 U546 ( .A1(n191), .A2(n137), .ZN(shiftedA_20__29_) );
  NOR2_X1 U547 ( .A1(n229), .A2(n100), .ZN(shiftedA_8__30_) );
  NOR2_X1 U548 ( .A1(n203), .A2(n128), .ZN(shiftedA_17__30_) );
  NOR2_X1 U549 ( .A1(n194), .A2(n137), .ZN(shiftedA_20__30_) );
  NOR2_X1 U550 ( .A1(n232), .A2(n100), .ZN(shiftedA_8__31_) );
  NOR2_X1 U551 ( .A1(n206), .A2(n128), .ZN(shiftedA_17__31_) );
  NOR2_X1 U552 ( .A1(n197), .A2(n137), .ZN(shiftedA_20__31_) );
  NOR2_X1 U553 ( .A1(n235), .A2(n100), .ZN(shiftedA_8__32_) );
  NOR2_X1 U554 ( .A1(n209), .A2(n128), .ZN(shiftedA_17__32_) );
  NOR2_X1 U555 ( .A1(n191), .A2(n146), .ZN(shiftedA_23__32_) );
  NOR2_X1 U556 ( .A1(n200), .A2(n137), .ZN(shiftedA_20__32_) );
  NOR2_X1 U557 ( .A1(n212), .A2(n128), .ZN(shiftedA_17__33_) );
  NOR2_X1 U558 ( .A1(n194), .A2(n146), .ZN(shiftedA_23__33_) );
  NOR2_X1 U559 ( .A1(n203), .A2(n137), .ZN(shiftedA_20__33_) );
  NOR2_X1 U560 ( .A1(n215), .A2(n128), .ZN(shiftedA_17__34_) );
  NOR2_X1 U561 ( .A1(n197), .A2(n146), .ZN(shiftedA_23__34_) );
  NOR2_X1 U562 ( .A1(n206), .A2(n137), .ZN(shiftedA_20__34_) );
  NOR2_X1 U563 ( .A1(n218), .A2(n128), .ZN(shiftedA_17__35_) );
  NOR2_X1 U564 ( .A1(n200), .A2(n146), .ZN(shiftedA_23__35_) );
  NOR2_X1 U565 ( .A1(n209), .A2(n137), .ZN(shiftedA_20__35_) );
  NOR2_X1 U566 ( .A1(n191), .A2(n155), .ZN(shiftedA_26__35_) );
  NOR2_X1 U567 ( .A1(n221), .A2(n127), .ZN(shiftedA_17__36_) );
  NOR2_X1 U568 ( .A1(n203), .A2(n146), .ZN(shiftedA_23__36_) );
  NOR2_X1 U569 ( .A1(n212), .A2(n137), .ZN(shiftedA_20__36_) );
  NOR2_X1 U570 ( .A1(n194), .A2(n155), .ZN(shiftedA_26__36_) );
  NOR2_X1 U571 ( .A1(n188), .A2(n164), .ZN(shiftedA_29__37_) );
  NOR2_X1 U572 ( .A1(n224), .A2(n127), .ZN(shiftedA_17__37_) );
  NOR2_X1 U573 ( .A1(n206), .A2(n146), .ZN(shiftedA_23__37_) );
  NOR2_X1 U574 ( .A1(n215), .A2(n137), .ZN(shiftedA_20__37_) );
  NOR2_X1 U575 ( .A1(n190), .A2(n164), .ZN(shiftedA_29__38_) );
  NOR2_X1 U576 ( .A1(n197), .A2(n155), .ZN(shiftedA_26__37_) );
  NOR2_X1 U577 ( .A1(n227), .A2(n127), .ZN(shiftedA_17__38_) );
  NOR2_X1 U578 ( .A1(n209), .A2(n146), .ZN(shiftedA_23__38_) );
  NOR2_X1 U579 ( .A1(n218), .A2(n137), .ZN(shiftedA_20__38_) );
  NOR2_X1 U580 ( .A1(n200), .A2(n155), .ZN(shiftedA_26__38_) );
  NOR2_X1 U581 ( .A1(n193), .A2(n164), .ZN(shiftedA_29__39_) );
  NOR2_X1 U582 ( .A1(n230), .A2(n127), .ZN(shiftedA_17__39_) );
  NOR2_X1 U583 ( .A1(n212), .A2(n146), .ZN(shiftedA_23__39_) );
  NOR2_X1 U584 ( .A1(n221), .A2(n136), .ZN(shiftedA_20__39_) );
  NOR2_X1 U585 ( .A1(n196), .A2(n164), .ZN(shiftedA_29__40_) );
  NOR2_X1 U586 ( .A1(n203), .A2(n155), .ZN(shiftedA_26__39_) );
  NOR2_X1 U587 ( .A1(n233), .A2(n127), .ZN(shiftedA_17__40_) );
  NOR2_X1 U588 ( .A1(n215), .A2(n146), .ZN(shiftedA_23__40_) );
  NOR2_X1 U589 ( .A1(n224), .A2(n136), .ZN(shiftedA_20__40_) );
  NOR2_X1 U590 ( .A1(n199), .A2(n164), .ZN(shiftedA_29__41_) );
  NOR2_X1 U591 ( .A1(n187), .A2(n137), .ZN(shiftedA_20__28_) );
  NOR2_X1 U592 ( .A1(n238), .A2(n91), .ZN(shiftedA_5__30_) );
  NOR2_X1 U593 ( .A1(n188), .A2(n146), .ZN(shiftedA_23__31_) );
  NOR2_X1 U594 ( .A1(n238), .A2(n100), .ZN(shiftedA_8__33_) );
  NOR2_X1 U595 ( .A1(n188), .A2(n155), .ZN(shiftedA_26__34_) );
  NOR2_X1 U596 ( .A1(n247), .A2(n84), .ZN(shiftedA_2__30_) );
  NOR2_X1 U597 ( .A1(n250), .A2(n84), .ZN(shiftedA_2__31_) );
  NOR2_X1 U598 ( .A1(n241), .A2(n91), .ZN(shiftedA_5__31_) );
  NOR2_X1 U599 ( .A1(n253), .A2(n84), .ZN(shiftedA_2__32_) );
  NOR2_X1 U600 ( .A1(n244), .A2(n91), .ZN(shiftedA_5__32_) );
  NOR2_X1 U601 ( .A1(n247), .A2(n91), .ZN(shiftedA_5__33_) );
  NOR2_X1 U602 ( .A1(n250), .A2(n91), .ZN(shiftedA_5__34_) );
  NOR2_X1 U603 ( .A1(n241), .A2(n100), .ZN(shiftedA_8__34_) );
  NOR2_X1 U604 ( .A1(n253), .A2(n91), .ZN(shiftedA_5__35_) );
  NOR2_X1 U605 ( .A1(n244), .A2(n100), .ZN(shiftedA_8__35_) );
  NOR2_X1 U606 ( .A1(n247), .A2(n100), .ZN(shiftedA_8__36_) );
  NOR2_X1 U607 ( .A1(n250), .A2(n100), .ZN(shiftedA_8__37_) );
  NOR2_X1 U608 ( .A1(n253), .A2(n100), .ZN(shiftedA_8__38_) );
  NOR2_X1 U609 ( .A1(n185), .A2(n146), .ZN(shiftedA_23__30_) );
  NOR2_X1 U610 ( .A1(n185), .A2(n155), .ZN(shiftedA_26__33_) );
  NOR2_X1 U611 ( .A1(n232), .A2(n94), .ZN(shiftedA_6__29_) );
  NOR2_X1 U612 ( .A1(n197), .A2(n131), .ZN(shiftedA_18__29_) );
  NOR2_X1 U613 ( .A1(n235), .A2(n94), .ZN(shiftedA_6__30_) );
  NOR2_X1 U614 ( .A1(n191), .A2(n140), .ZN(shiftedA_21__30_) );
  NOR2_X1 U615 ( .A1(n200), .A2(n131), .ZN(shiftedA_18__30_) );
  NOR2_X1 U616 ( .A1(n103), .A2(n229), .ZN(shiftedA_9__31_) );
  NOR2_X1 U617 ( .A1(n194), .A2(n140), .ZN(shiftedA_21__31_) );
  NOR2_X1 U618 ( .A1(n203), .A2(n131), .ZN(shiftedA_18__31_) );
  NOR2_X1 U619 ( .A1(n103), .A2(n232), .ZN(shiftedA_9__32_) );
  NOR2_X1 U620 ( .A1(n197), .A2(n140), .ZN(shiftedA_21__32_) );
  NOR2_X1 U621 ( .A1(n206), .A2(n131), .ZN(shiftedA_18__32_) );
  NOR2_X1 U622 ( .A1(n103), .A2(n235), .ZN(shiftedA_9__33_) );
  NOR2_X1 U623 ( .A1(n200), .A2(n140), .ZN(shiftedA_21__33_) );
  NOR2_X1 U624 ( .A1(n209), .A2(n131), .ZN(shiftedA_18__33_) );
  NOR2_X1 U625 ( .A1(n103), .A2(n238), .ZN(shiftedA_9__34_) );
  NOR2_X1 U626 ( .A1(n191), .A2(n149), .ZN(shiftedA_24__33_) );
  NOR2_X1 U627 ( .A1(n203), .A2(n140), .ZN(shiftedA_21__34_) );
  NOR2_X1 U628 ( .A1(n212), .A2(n131), .ZN(shiftedA_18__34_) );
  NOR2_X1 U629 ( .A1(n103), .A2(n241), .ZN(shiftedA_9__35_) );
  NOR2_X1 U630 ( .A1(n188), .A2(n158), .ZN(shiftedA_27__35_) );
  NOR2_X1 U631 ( .A1(n194), .A2(n149), .ZN(shiftedA_24__34_) );
  NOR2_X1 U632 ( .A1(n206), .A2(n140), .ZN(shiftedA_21__35_) );
  NOR2_X1 U633 ( .A1(n215), .A2(n131), .ZN(shiftedA_18__35_) );
  NOR2_X1 U634 ( .A1(n190), .A2(n158), .ZN(shiftedA_27__36_) );
  NOR2_X1 U635 ( .A1(n103), .A2(n244), .ZN(shiftedA_9__36_) );
  NOR2_X1 U636 ( .A1(n197), .A2(n149), .ZN(shiftedA_24__35_) );
  NOR2_X1 U637 ( .A1(n209), .A2(n140), .ZN(shiftedA_21__36_) );
  NOR2_X1 U638 ( .A1(n218), .A2(n131), .ZN(shiftedA_18__36_) );
  NOR2_X1 U639 ( .A1(n200), .A2(n149), .ZN(shiftedA_24__36_) );
  NOR2_X1 U640 ( .A1(n103), .A2(n247), .ZN(shiftedA_9__37_) );
  NOR2_X1 U641 ( .A1(n193), .A2(n158), .ZN(shiftedA_27__37_) );
  NOR2_X1 U642 ( .A1(n212), .A2(n140), .ZN(shiftedA_21__37_) );
  NOR2_X1 U643 ( .A1(n221), .A2(n130), .ZN(shiftedA_18__37_) );
  NOR2_X1 U644 ( .A1(n187), .A2(n167), .ZN(shiftedA_30__38_) );
  NOR2_X1 U645 ( .A1(n196), .A2(n158), .ZN(shiftedA_27__38_) );
  NOR2_X1 U646 ( .A1(n103), .A2(n250), .ZN(shiftedA_9__38_) );
  NOR2_X1 U647 ( .A1(n203), .A2(n149), .ZN(shiftedA_24__37_) );
  NOR2_X1 U648 ( .A1(n215), .A2(n140), .ZN(shiftedA_21__38_) );
  NOR2_X1 U649 ( .A1(n224), .A2(n130), .ZN(shiftedA_18__38_) );
  NOR2_X1 U650 ( .A1(n206), .A2(n149), .ZN(shiftedA_24__38_) );
  NOR2_X1 U651 ( .A1(n103), .A2(n253), .ZN(shiftedA_9__39_) );
  NOR2_X1 U652 ( .A1(n190), .A2(n167), .ZN(shiftedA_30__39_) );
  NOR2_X1 U653 ( .A1(n199), .A2(n158), .ZN(shiftedA_27__39_) );
  NOR2_X1 U654 ( .A1(n218), .A2(n140), .ZN(shiftedA_21__39_) );
  NOR2_X1 U655 ( .A1(n227), .A2(n130), .ZN(shiftedA_18__39_) );
  NOR2_X1 U656 ( .A1(n193), .A2(n167), .ZN(shiftedA_30__40_) );
  NOR2_X1 U657 ( .A1(n202), .A2(n158), .ZN(shiftedA_27__40_) );
  NOR2_X1 U658 ( .A1(n209), .A2(n149), .ZN(shiftedA_24__39_) );
  NOR2_X1 U659 ( .A1(n221), .A2(n139), .ZN(shiftedA_21__40_) );
  NOR2_X1 U660 ( .A1(n230), .A2(n130), .ZN(shiftedA_18__40_) );
  NOR2_X1 U661 ( .A1(n196), .A2(n167), .ZN(shiftedA_30__41_) );
  NOR2_X1 U662 ( .A1(n205), .A2(n158), .ZN(shiftedA_27__41_) );
  NOR2_X1 U663 ( .A1(n212), .A2(n149), .ZN(shiftedA_24__40_) );
  NOR2_X1 U664 ( .A1(n224), .A2(n139), .ZN(shiftedA_21__41_) );
  NOR2_X1 U665 ( .A1(n233), .A2(n130), .ZN(shiftedA_18__41_) );
  NOR2_X1 U666 ( .A1(n199), .A2(n167), .ZN(shiftedA_30__42_) );
  NOR2_X1 U667 ( .A1(n208), .A2(n158), .ZN(shiftedA_27__42_) );
  NOR2_X1 U668 ( .A1(n238), .A2(n94), .ZN(shiftedA_6__31_) );
  NOR2_X1 U669 ( .A1(n187), .A2(n149), .ZN(shiftedA_24__32_) );
  NOR2_X1 U670 ( .A1(n241), .A2(n94), .ZN(shiftedA_6__32_) );
  NOR2_X1 U671 ( .A1(n244), .A2(n94), .ZN(shiftedA_6__33_) );
  NOR2_X1 U672 ( .A1(n247), .A2(n94), .ZN(shiftedA_6__34_) );
  NOR2_X1 U673 ( .A1(n250), .A2(n94), .ZN(shiftedA_6__35_) );
  NOR2_X1 U674 ( .A1(n253), .A2(n94), .ZN(shiftedA_6__36_) );
  NOR2_X1 U675 ( .A1(n185), .A2(n158), .ZN(shiftedA_27__34_) );
  NOR2_X1 U676 ( .A1(n182), .A2(n162), .ZN(shiftedA_28__34_) );
  NOR2_X1 U677 ( .A1(n229), .A2(n97), .ZN(shiftedA_7__29_) );
  NOR2_X1 U678 ( .A1(n203), .A2(n125), .ZN(shiftedA_16__29_) );
  NOR2_X1 U679 ( .A1(n194), .A2(n134), .ZN(shiftedA_19__29_) );
  NOR2_X1 U680 ( .A1(n232), .A2(n97), .ZN(shiftedA_7__30_) );
  NOR2_X1 U681 ( .A1(n206), .A2(n125), .ZN(shiftedA_16__30_) );
  NOR2_X1 U682 ( .A1(n197), .A2(n134), .ZN(shiftedA_19__30_) );
  NOR2_X1 U683 ( .A1(n235), .A2(n97), .ZN(shiftedA_7__31_) );
  NOR2_X1 U684 ( .A1(n209), .A2(n125), .ZN(shiftedA_16__31_) );
  NOR2_X1 U685 ( .A1(n191), .A2(n143), .ZN(shiftedA_22__31_) );
  NOR2_X1 U686 ( .A1(n200), .A2(n134), .ZN(shiftedA_19__31_) );
  NOR2_X1 U687 ( .A1(n212), .A2(n125), .ZN(shiftedA_16__32_) );
  NOR2_X1 U688 ( .A1(n194), .A2(n143), .ZN(shiftedA_22__32_) );
  NOR2_X1 U689 ( .A1(n203), .A2(n134), .ZN(shiftedA_19__32_) );
  NOR2_X1 U690 ( .A1(n215), .A2(n125), .ZN(shiftedA_16__33_) );
  NOR2_X1 U691 ( .A1(n197), .A2(n143), .ZN(shiftedA_22__33_) );
  NOR2_X1 U692 ( .A1(n206), .A2(n134), .ZN(shiftedA_19__33_) );
  NOR2_X1 U693 ( .A1(n218), .A2(n125), .ZN(shiftedA_16__34_) );
  NOR2_X1 U694 ( .A1(n200), .A2(n143), .ZN(shiftedA_22__34_) );
  NOR2_X1 U695 ( .A1(n209), .A2(n134), .ZN(shiftedA_19__34_) );
  NOR2_X1 U696 ( .A1(n191), .A2(n152), .ZN(shiftedA_25__34_) );
  NOR2_X1 U697 ( .A1(n221), .A2(n124), .ZN(shiftedA_16__35_) );
  NOR2_X1 U698 ( .A1(n203), .A2(n143), .ZN(shiftedA_22__35_) );
  NOR2_X1 U699 ( .A1(n212), .A2(n134), .ZN(shiftedA_19__35_) );
  NOR2_X1 U700 ( .A1(n187), .A2(n161), .ZN(shiftedA_28__36_) );
  NOR2_X1 U701 ( .A1(n194), .A2(n152), .ZN(shiftedA_25__35_) );
  NOR2_X1 U702 ( .A1(n224), .A2(n124), .ZN(shiftedA_16__36_) );
  NOR2_X1 U703 ( .A1(n206), .A2(n143), .ZN(shiftedA_22__36_) );
  NOR2_X1 U704 ( .A1(n215), .A2(n134), .ZN(shiftedA_19__36_) );
  NOR2_X1 U705 ( .A1(n197), .A2(n152), .ZN(shiftedA_25__36_) );
  NOR2_X1 U706 ( .A1(n190), .A2(n161), .ZN(shiftedA_28__37_) );
  NOR2_X1 U707 ( .A1(n227), .A2(n124), .ZN(shiftedA_16__37_) );
  NOR2_X1 U708 ( .A1(n209), .A2(n143), .ZN(shiftedA_22__37_) );
  NOR2_X1 U709 ( .A1(n218), .A2(n134), .ZN(shiftedA_19__37_) );
  NOR2_X1 U710 ( .A1(n193), .A2(n161), .ZN(shiftedA_28__38_) );
  NOR2_X1 U711 ( .A1(n200), .A2(n152), .ZN(shiftedA_25__37_) );
  NOR2_X1 U712 ( .A1(n230), .A2(n124), .ZN(shiftedA_16__38_) );
  NOR2_X1 U713 ( .A1(n212), .A2(n143), .ZN(shiftedA_22__38_) );
  NOR2_X1 U714 ( .A1(n221), .A2(n133), .ZN(shiftedA_19__38_) );
  NOR2_X1 U715 ( .A1(n203), .A2(n152), .ZN(shiftedA_25__38_) );
  NOR2_X1 U716 ( .A1(n196), .A2(n161), .ZN(shiftedA_28__39_) );
  NOR2_X1 U717 ( .A1(n233), .A2(n124), .ZN(shiftedA_16__39_) );
  NOR2_X1 U718 ( .A1(n215), .A2(n143), .ZN(shiftedA_22__39_) );
  NOR2_X1 U719 ( .A1(n224), .A2(n133), .ZN(shiftedA_19__39_) );
  NOR2_X1 U720 ( .A1(n199), .A2(n161), .ZN(shiftedA_28__40_) );
  NOR2_X1 U721 ( .A1(n206), .A2(n152), .ZN(shiftedA_25__39_) );
  NOR2_X1 U722 ( .A1(n236), .A2(n124), .ZN(shiftedA_16__40_) );
  NOR2_X1 U723 ( .A1(n218), .A2(n143), .ZN(shiftedA_22__40_) );
  NOR2_X1 U724 ( .A1(n227), .A2(n133), .ZN(shiftedA_19__40_) );
  NOR2_X1 U725 ( .A1(n202), .A2(n161), .ZN(shiftedA_28__41_) );
  NOR2_X1 U726 ( .A1(n209), .A2(n152), .ZN(shiftedA_25__40_) );
  NOR2_X1 U727 ( .A1(n239), .A2(n124), .ZN(shiftedA_16__41_) );
  NOR2_X1 U728 ( .A1(n221), .A2(n142), .ZN(shiftedA_22__41_) );
  NOR2_X1 U729 ( .A1(n230), .A2(n133), .ZN(shiftedA_19__41_) );
  NOR2_X1 U730 ( .A1(n205), .A2(n161), .ZN(shiftedA_28__42_) );
  NOR2_X1 U731 ( .A1(n188), .A2(n143), .ZN(shiftedA_22__30_) );
  NOR2_X1 U732 ( .A1(n238), .A2(n97), .ZN(shiftedA_7__32_) );
  NOR2_X1 U733 ( .A1(n188), .A2(n152), .ZN(shiftedA_25__33_) );
  NOR2_X1 U734 ( .A1(n241), .A2(n97), .ZN(shiftedA_7__33_) );
  NOR2_X1 U735 ( .A1(n244), .A2(n97), .ZN(shiftedA_7__34_) );
  NOR2_X1 U736 ( .A1(n247), .A2(n97), .ZN(shiftedA_7__35_) );
  NOR2_X1 U737 ( .A1(n250), .A2(n97), .ZN(shiftedA_7__36_) );
  NOR2_X1 U738 ( .A1(n253), .A2(n97), .ZN(shiftedA_7__37_) );
  NOR2_X1 U739 ( .A1(n249), .A2(n118), .ZN(shiftedA_14__42_) );
  NOR2_X1 U740 ( .A1(n252), .A2(n118), .ZN(shiftedA_14__43_) );
  NOR2_X1 U741 ( .A1(n255), .A2(n118), .ZN(shiftedA_14__44_) );
  NOR2_X1 U742 ( .A1(n246), .A2(n121), .ZN(shiftedA_15__42_) );
  NOR2_X1 U743 ( .A1(n249), .A2(n121), .ZN(shiftedA_15__43_) );
  NOR2_X1 U744 ( .A1(n252), .A2(n121), .ZN(shiftedA_15__44_) );
  NOR2_X1 U745 ( .A1(n255), .A2(n121), .ZN(shiftedA_15__45_) );
  NOR2_X1 U746 ( .A1(n255), .A2(n115), .ZN(shiftedA_13__43_) );
  NOR2_X1 U747 ( .A1(n206), .A2(n155), .ZN(shiftedA_26__40_) );
  NOR2_X1 U748 ( .A1(n236), .A2(n127), .ZN(shiftedA_17__41_) );
  NOR2_X1 U749 ( .A1(n218), .A2(n146), .ZN(shiftedA_23__41_) );
  NOR2_X1 U750 ( .A1(n227), .A2(n136), .ZN(shiftedA_20__41_) );
  NOR2_X1 U751 ( .A1(n202), .A2(n164), .ZN(shiftedA_29__42_) );
  NOR2_X1 U752 ( .A1(n209), .A2(n155), .ZN(shiftedA_26__41_) );
  NOR2_X1 U753 ( .A1(n239), .A2(n127), .ZN(shiftedA_17__42_) );
  NOR2_X1 U754 ( .A1(n221), .A2(n145), .ZN(shiftedA_23__42_) );
  NOR2_X1 U755 ( .A1(n230), .A2(n136), .ZN(shiftedA_20__42_) );
  NOR2_X1 U756 ( .A1(n205), .A2(n164), .ZN(shiftedA_29__43_) );
  NOR2_X1 U757 ( .A1(n212), .A2(n155), .ZN(shiftedA_26__42_) );
  NOR2_X1 U758 ( .A1(n242), .A2(n127), .ZN(shiftedA_17__43_) );
  NOR2_X1 U759 ( .A1(n224), .A2(n145), .ZN(shiftedA_23__43_) );
  NOR2_X1 U760 ( .A1(n233), .A2(n136), .ZN(shiftedA_20__43_) );
  NOR2_X1 U761 ( .A1(n208), .A2(n164), .ZN(shiftedA_29__44_) );
  NOR2_X1 U762 ( .A1(n215), .A2(n155), .ZN(shiftedA_26__43_) );
  NOR2_X1 U763 ( .A1(n227), .A2(n145), .ZN(shiftedA_23__44_) );
  NOR2_X1 U764 ( .A1(n236), .A2(n136), .ZN(shiftedA_20__44_) );
  NOR2_X1 U765 ( .A1(n211), .A2(n164), .ZN(shiftedA_29__45_) );
  NOR2_X1 U766 ( .A1(n218), .A2(n155), .ZN(shiftedA_26__44_) );
  NOR2_X1 U767 ( .A1(n230), .A2(n145), .ZN(shiftedA_23__45_) );
  NOR2_X1 U768 ( .A1(n239), .A2(n136), .ZN(shiftedA_20__45_) );
  NOR2_X1 U769 ( .A1(n214), .A2(n164), .ZN(shiftedA_29__46_) );
  NOR2_X1 U770 ( .A1(n221), .A2(n154), .ZN(shiftedA_26__45_) );
  NOR2_X1 U771 ( .A1(n233), .A2(n145), .ZN(shiftedA_23__46_) );
  NOR2_X1 U772 ( .A1(n242), .A2(n136), .ZN(shiftedA_20__46_) );
  NOR2_X1 U773 ( .A1(n217), .A2(n164), .ZN(shiftedA_29__47_) );
  NOR2_X1 U774 ( .A1(n224), .A2(n154), .ZN(shiftedA_26__46_) );
  NOR2_X1 U775 ( .A1(n236), .A2(n145), .ZN(shiftedA_23__47_) );
  NOR2_X1 U776 ( .A1(n220), .A2(n163), .ZN(shiftedA_29__48_) );
  NOR2_X1 U777 ( .A1(n227), .A2(n154), .ZN(shiftedA_26__47_) );
  NOR2_X1 U778 ( .A1(n239), .A2(n145), .ZN(shiftedA_23__48_) );
  NOR2_X1 U779 ( .A1(n223), .A2(n163), .ZN(shiftedA_29__49_) );
  NOR2_X1 U780 ( .A1(n230), .A2(n154), .ZN(shiftedA_26__48_) );
  NOR2_X1 U781 ( .A1(n242), .A2(n145), .ZN(shiftedA_23__49_) );
  NOR2_X1 U782 ( .A1(n226), .A2(n163), .ZN(shiftedA_29__50_) );
  NOR2_X1 U783 ( .A1(n233), .A2(n154), .ZN(shiftedA_26__49_) );
  NOR2_X1 U784 ( .A1(n229), .A2(n163), .ZN(shiftedA_29__51_) );
  NOR2_X1 U785 ( .A1(n236), .A2(n154), .ZN(shiftedA_26__50_) );
  NOR2_X1 U786 ( .A1(n239), .A2(n154), .ZN(shiftedA_26__51_) );
  NOR2_X1 U787 ( .A1(n232), .A2(n163), .ZN(shiftedA_29__52_) );
  NOR2_X1 U788 ( .A1(n235), .A2(n163), .ZN(shiftedA_29__53_) );
  NOR2_X1 U789 ( .A1(n242), .A2(n154), .ZN(shiftedA_26__52_) );
  NOR2_X1 U790 ( .A1(n245), .A2(n127), .ZN(shiftedA_17__44_) );
  NOR2_X1 U791 ( .A1(n248), .A2(n127), .ZN(shiftedA_17__45_) );
  NOR2_X1 U792 ( .A1(n251), .A2(n127), .ZN(shiftedA_17__46_) );
  NOR2_X1 U793 ( .A1(n254), .A2(n127), .ZN(shiftedA_17__47_) );
  NOR2_X1 U794 ( .A1(n245), .A2(n136), .ZN(shiftedA_20__47_) );
  NOR2_X1 U795 ( .A1(n248), .A2(n136), .ZN(shiftedA_20__48_) );
  NOR2_X1 U796 ( .A1(n251), .A2(n136), .ZN(shiftedA_20__49_) );
  NOR2_X1 U797 ( .A1(n254), .A2(n136), .ZN(shiftedA_20__50_) );
  NOR2_X1 U798 ( .A1(n245), .A2(n145), .ZN(shiftedA_23__50_) );
  NOR2_X1 U799 ( .A1(n248), .A2(n145), .ZN(shiftedA_23__51_) );
  NOR2_X1 U800 ( .A1(n251), .A2(n145), .ZN(shiftedA_23__52_) );
  NOR2_X1 U801 ( .A1(n254), .A2(n145), .ZN(shiftedA_23__53_) );
  NOR2_X1 U802 ( .A1(n238), .A2(n163), .ZN(shiftedA_29__54_) );
  NOR2_X1 U803 ( .A1(n215), .A2(n149), .ZN(shiftedA_24__41_) );
  NOR2_X1 U804 ( .A1(n227), .A2(n139), .ZN(shiftedA_21__42_) );
  NOR2_X1 U805 ( .A1(n236), .A2(n130), .ZN(shiftedA_18__42_) );
  NOR2_X1 U806 ( .A1(n202), .A2(n167), .ZN(shiftedA_30__43_) );
  NOR2_X1 U807 ( .A1(n211), .A2(n158), .ZN(shiftedA_27__43_) );
  NOR2_X1 U808 ( .A1(n218), .A2(n149), .ZN(shiftedA_24__42_) );
  NOR2_X1 U809 ( .A1(n230), .A2(n139), .ZN(shiftedA_21__43_) );
  NOR2_X1 U810 ( .A1(n239), .A2(n130), .ZN(shiftedA_18__43_) );
  NOR2_X1 U811 ( .A1(n205), .A2(n167), .ZN(shiftedA_30__44_) );
  NOR2_X1 U812 ( .A1(n214), .A2(n158), .ZN(shiftedA_27__44_) );
  NOR2_X1 U813 ( .A1(n221), .A2(n148), .ZN(shiftedA_24__43_) );
  NOR2_X1 U814 ( .A1(n233), .A2(n139), .ZN(shiftedA_21__44_) );
  NOR2_X1 U815 ( .A1(n242), .A2(n130), .ZN(shiftedA_18__44_) );
  NOR2_X1 U816 ( .A1(n208), .A2(n167), .ZN(shiftedA_30__45_) );
  NOR2_X1 U817 ( .A1(n217), .A2(n158), .ZN(shiftedA_27__45_) );
  NOR2_X1 U818 ( .A1(n224), .A2(n148), .ZN(shiftedA_24__44_) );
  NOR2_X1 U819 ( .A1(n236), .A2(n139), .ZN(shiftedA_21__45_) );
  NOR2_X1 U820 ( .A1(n211), .A2(n167), .ZN(shiftedA_30__46_) );
  NOR2_X1 U821 ( .A1(n220), .A2(n157), .ZN(shiftedA_27__46_) );
  NOR2_X1 U822 ( .A1(n227), .A2(n148), .ZN(shiftedA_24__45_) );
  NOR2_X1 U823 ( .A1(n239), .A2(n139), .ZN(shiftedA_21__46_) );
  NOR2_X1 U824 ( .A1(n214), .A2(n167), .ZN(shiftedA_30__47_) );
  NOR2_X1 U825 ( .A1(n223), .A2(n157), .ZN(shiftedA_27__47_) );
  NOR2_X1 U826 ( .A1(n230), .A2(n148), .ZN(shiftedA_24__46_) );
  NOR2_X1 U827 ( .A1(n242), .A2(n139), .ZN(shiftedA_21__47_) );
  NOR2_X1 U828 ( .A1(n217), .A2(n167), .ZN(shiftedA_30__48_) );
  NOR2_X1 U829 ( .A1(n226), .A2(n157), .ZN(shiftedA_27__48_) );
  NOR2_X1 U830 ( .A1(n233), .A2(n148), .ZN(shiftedA_24__47_) );
  NOR2_X1 U831 ( .A1(n220), .A2(n166), .ZN(shiftedA_30__49_) );
  NOR2_X1 U832 ( .A1(n229), .A2(n157), .ZN(shiftedA_27__49_) );
  NOR2_X1 U833 ( .A1(n236), .A2(n148), .ZN(shiftedA_24__48_) );
  NOR2_X1 U834 ( .A1(n223), .A2(n166), .ZN(shiftedA_30__50_) );
  NOR2_X1 U835 ( .A1(n232), .A2(n157), .ZN(shiftedA_27__50_) );
  NOR2_X1 U836 ( .A1(n239), .A2(n148), .ZN(shiftedA_24__49_) );
  NOR2_X1 U837 ( .A1(n226), .A2(n166), .ZN(shiftedA_30__51_) );
  NOR2_X1 U838 ( .A1(n235), .A2(n157), .ZN(shiftedA_27__51_) );
  NOR2_X1 U839 ( .A1(n242), .A2(n148), .ZN(shiftedA_24__50_) );
  NOR2_X1 U840 ( .A1(n229), .A2(n166), .ZN(shiftedA_30__52_) );
  NOR2_X1 U841 ( .A1(n232), .A2(n166), .ZN(shiftedA_30__53_) );
  NOR2_X1 U842 ( .A1(n235), .A2(n166), .ZN(shiftedA_30__54_) );
  NOR2_X1 U843 ( .A1(n245), .A2(n130), .ZN(shiftedA_18__45_) );
  NOR2_X1 U844 ( .A1(n248), .A2(n130), .ZN(shiftedA_18__46_) );
  NOR2_X1 U845 ( .A1(n251), .A2(n130), .ZN(shiftedA_18__47_) );
  NOR2_X1 U846 ( .A1(n245), .A2(n139), .ZN(shiftedA_21__48_) );
  NOR2_X1 U847 ( .A1(n254), .A2(n130), .ZN(shiftedA_18__48_) );
  NOR2_X1 U848 ( .A1(n248), .A2(n139), .ZN(shiftedA_21__49_) );
  NOR2_X1 U849 ( .A1(n251), .A2(n139), .ZN(shiftedA_21__50_) );
  NOR2_X1 U850 ( .A1(n254), .A2(n139), .ZN(shiftedA_21__51_) );
  NOR2_X1 U851 ( .A1(n245), .A2(n148), .ZN(shiftedA_24__51_) );
  NOR2_X1 U852 ( .A1(n238), .A2(n157), .ZN(shiftedA_27__52_) );
  NOR2_X1 U853 ( .A1(n248), .A2(n148), .ZN(shiftedA_24__52_) );
  NOR2_X1 U854 ( .A1(n251), .A2(n148), .ZN(shiftedA_24__53_) );
  NOR2_X1 U855 ( .A1(n238), .A2(n166), .ZN(shiftedA_30__55_) );
  NOR2_X1 U856 ( .A1(n241), .A2(n157), .ZN(shiftedA_27__53_) );
  NOR2_X1 U857 ( .A1(n244), .A2(n157), .ZN(shiftedA_27__54_) );
  NOR2_X1 U858 ( .A1(n247), .A2(n157), .ZN(shiftedA_27__55_) );
  NOR2_X1 U859 ( .A1(n212), .A2(n152), .ZN(shiftedA_25__41_) );
  NOR2_X1 U860 ( .A1(n242), .A2(n124), .ZN(shiftedA_16__42_) );
  NOR2_X1 U861 ( .A1(n224), .A2(n142), .ZN(shiftedA_22__42_) );
  NOR2_X1 U862 ( .A1(n233), .A2(n133), .ZN(shiftedA_19__42_) );
  NOR2_X1 U863 ( .A1(n208), .A2(n161), .ZN(shiftedA_28__43_) );
  NOR2_X1 U864 ( .A1(n215), .A2(n152), .ZN(shiftedA_25__42_) );
  NOR2_X1 U865 ( .A1(n227), .A2(n142), .ZN(shiftedA_22__43_) );
  NOR2_X1 U866 ( .A1(n236), .A2(n133), .ZN(shiftedA_19__43_) );
  NOR2_X1 U867 ( .A1(n211), .A2(n161), .ZN(shiftedA_28__44_) );
  NOR2_X1 U868 ( .A1(n218), .A2(n152), .ZN(shiftedA_25__43_) );
  NOR2_X1 U869 ( .A1(n230), .A2(n142), .ZN(shiftedA_22__44_) );
  NOR2_X1 U870 ( .A1(n239), .A2(n133), .ZN(shiftedA_19__44_) );
  NOR2_X1 U871 ( .A1(n214), .A2(n161), .ZN(shiftedA_28__45_) );
  NOR2_X1 U872 ( .A1(n221), .A2(n151), .ZN(shiftedA_25__44_) );
  NOR2_X1 U873 ( .A1(n233), .A2(n142), .ZN(shiftedA_22__45_) );
  NOR2_X1 U874 ( .A1(n242), .A2(n133), .ZN(shiftedA_19__45_) );
  NOR2_X1 U875 ( .A1(n217), .A2(n161), .ZN(shiftedA_28__46_) );
  NOR2_X1 U876 ( .A1(n224), .A2(n151), .ZN(shiftedA_25__45_) );
  NOR2_X1 U877 ( .A1(n236), .A2(n142), .ZN(shiftedA_22__46_) );
  NOR2_X1 U878 ( .A1(n220), .A2(n160), .ZN(shiftedA_28__47_) );
  NOR2_X1 U879 ( .A1(n227), .A2(n151), .ZN(shiftedA_25__46_) );
  NOR2_X1 U880 ( .A1(n239), .A2(n142), .ZN(shiftedA_22__47_) );
  NOR2_X1 U881 ( .A1(n223), .A2(n160), .ZN(shiftedA_28__48_) );
  NOR2_X1 U882 ( .A1(n230), .A2(n151), .ZN(shiftedA_25__47_) );
  NOR2_X1 U883 ( .A1(n242), .A2(n142), .ZN(shiftedA_22__48_) );
  NOR2_X1 U884 ( .A1(n226), .A2(n160), .ZN(shiftedA_28__49_) );
  NOR2_X1 U885 ( .A1(n233), .A2(n151), .ZN(shiftedA_25__48_) );
  NOR2_X1 U886 ( .A1(n229), .A2(n160), .ZN(shiftedA_28__50_) );
  NOR2_X1 U887 ( .A1(n236), .A2(n151), .ZN(shiftedA_25__49_) );
  NOR2_X1 U888 ( .A1(n232), .A2(n160), .ZN(shiftedA_28__51_) );
  NOR2_X1 U889 ( .A1(n239), .A2(n151), .ZN(shiftedA_25__50_) );
  NOR2_X1 U890 ( .A1(n242), .A2(n151), .ZN(shiftedA_25__51_) );
  NOR2_X1 U891 ( .A1(n235), .A2(n160), .ZN(shiftedA_28__52_) );
  NOR2_X1 U892 ( .A1(n245), .A2(n124), .ZN(shiftedA_16__43_) );
  NOR2_X1 U893 ( .A1(n248), .A2(n124), .ZN(shiftedA_16__44_) );
  NOR2_X1 U894 ( .A1(n251), .A2(n124), .ZN(shiftedA_16__45_) );
  NOR2_X1 U895 ( .A1(n254), .A2(n124), .ZN(shiftedA_16__46_) );
  NOR2_X1 U896 ( .A1(n245), .A2(n133), .ZN(shiftedA_19__46_) );
  NOR2_X1 U897 ( .A1(n248), .A2(n133), .ZN(shiftedA_19__47_) );
  NOR2_X1 U898 ( .A1(n251), .A2(n133), .ZN(shiftedA_19__48_) );
  NOR2_X1 U899 ( .A1(n254), .A2(n133), .ZN(shiftedA_19__49_) );
  NOR2_X1 U900 ( .A1(n245), .A2(n142), .ZN(shiftedA_22__49_) );
  NOR2_X1 U901 ( .A1(n248), .A2(n142), .ZN(shiftedA_22__50_) );
  NOR2_X1 U902 ( .A1(n251), .A2(n142), .ZN(shiftedA_22__51_) );
  NOR2_X1 U903 ( .A1(n254), .A2(n142), .ZN(shiftedA_22__52_) );
  NOR2_X1 U904 ( .A1(n238), .A2(n160), .ZN(shiftedA_28__53_) );
  NOR2_X1 U905 ( .A1(n245), .A2(n151), .ZN(shiftedA_25__52_) );
  NOR2_X1 U906 ( .A1(n248), .A2(n151), .ZN(shiftedA_25__53_) );
  NOR2_X1 U907 ( .A1(n241), .A2(n160), .ZN(shiftedA_28__54_) );
  NOR2_X1 U908 ( .A1(n244), .A2(n160), .ZN(shiftedA_28__55_) );
  BUF_X1 U909 ( .A(shiftedA_56__63_), .Z(n324) );
  NOR2_X1 U910 ( .A1(n171), .A2(n81), .ZN(shiftedA_0__0_) );
  NOR2_X1 U911 ( .A1(n245), .A2(n154), .ZN(shiftedA_26__53_) );
  NOR2_X1 U912 ( .A1(n248), .A2(n154), .ZN(shiftedA_26__54_) );
  NOR2_X1 U913 ( .A1(n251), .A2(n154), .ZN(shiftedA_26__55_) );
  NOR2_X1 U914 ( .A1(n254), .A2(n154), .ZN(shiftedA_26__56_) );
  NOR2_X1 U915 ( .A1(n241), .A2(n163), .ZN(shiftedA_29__55_) );
  NOR2_X1 U916 ( .A1(n244), .A2(n163), .ZN(shiftedA_29__56_) );
  NOR2_X1 U917 ( .A1(n247), .A2(n163), .ZN(shiftedA_29__57_) );
  NOR2_X1 U918 ( .A1(n250), .A2(n163), .ZN(shiftedA_29__58_) );
  NOR2_X1 U919 ( .A1(n253), .A2(n163), .ZN(shiftedA_29__59_) );
  NOR2_X1 U920 ( .A1(n254), .A2(n148), .ZN(shiftedA_24__54_) );
  NOR2_X1 U921 ( .A1(n241), .A2(n166), .ZN(shiftedA_30__56_) );
  NOR2_X1 U922 ( .A1(n250), .A2(n157), .ZN(shiftedA_27__56_) );
  NOR2_X1 U923 ( .A1(n244), .A2(n166), .ZN(shiftedA_30__57_) );
  NOR2_X1 U924 ( .A1(n253), .A2(n157), .ZN(shiftedA_27__57_) );
  NOR2_X1 U925 ( .A1(n247), .A2(n166), .ZN(shiftedA_30__58_) );
  NOR2_X1 U926 ( .A1(n250), .A2(n166), .ZN(shiftedA_30__59_) );
  NOR2_X1 U927 ( .A1(n253), .A2(n166), .ZN(shiftedA_30__60_) );
  NOR2_X1 U928 ( .A1(n251), .A2(n151), .ZN(shiftedA_25__54_) );
  NOR2_X1 U929 ( .A1(n254), .A2(n151), .ZN(shiftedA_25__55_) );
  NOR2_X1 U930 ( .A1(n247), .A2(n160), .ZN(shiftedA_28__56_) );
  NOR2_X1 U931 ( .A1(n250), .A2(n160), .ZN(shiftedA_28__57_) );
  NOR2_X1 U932 ( .A1(n253), .A2(n160), .ZN(shiftedA_28__58_) );
  BUF_X2 U933 ( .A(shiftedA_0__63_), .Z(n346) );
  BUF_X2 U934 ( .A(n59), .Z(n87) );
  BUF_X1 U935 ( .A(n31), .Z(n171) );
  BUF_X1 U936 ( .A(n20), .Z(n198) );
  BUF_X1 U937 ( .A(n21), .Z(n195) );
  BUF_X1 U938 ( .A(n19), .Z(n201) );
  BUF_X1 U939 ( .A(n13), .Z(n219) );
  BUF_X1 U940 ( .A(n18), .Z(n204) );
  BUF_X1 U941 ( .A(n12), .Z(n222) );
  BUF_X1 U942 ( .A(n17), .Z(n207) );
  BUF_X1 U943 ( .A(n16), .Z(n210) );
  BUF_X1 U944 ( .A(n15), .Z(n213) );
  BUF_X1 U945 ( .A(n14), .Z(n216) );
  BUF_X1 U946 ( .A(n11), .Z(n225) );
  BUF_X1 U947 ( .A(n10), .Z(n228) );
  BUF_X1 U948 ( .A(n9), .Z(n231) );
  BUF_X1 U949 ( .A(n8), .Z(n234) );
  BUF_X1 U950 ( .A(n7), .Z(n237) );
  BUF_X1 U951 ( .A(n6), .Z(n240) );
  BUF_X1 U952 ( .A(n5), .Z(n243) );
  BUF_X1 U953 ( .A(n51), .Z(n111) );
  BUF_X1 U954 ( .A(n49), .Z(n117) );
  BUF_X1 U955 ( .A(n45), .Z(n129) );
  BUF_X1 U956 ( .A(n47), .Z(n123) );
  BUF_X1 U957 ( .A(n46), .Z(n126) );
  BUF_X1 U958 ( .A(n42), .Z(n138) );
  BUF_X1 U959 ( .A(n41), .Z(n141) );
  BUF_X1 U960 ( .A(n39), .Z(n147) );
  BUF_X1 U961 ( .A(n37), .Z(n153) );
  BUF_X1 U962 ( .A(n36), .Z(n156) );
  CLKBUF_X1 U963 ( .A(n24), .Z(n77) );
  BUF_X1 U964 ( .A(n4), .Z(n246) );
  BUF_X1 U965 ( .A(n3), .Z(n249) );
  BUF_X1 U966 ( .A(n2), .Z(n252) );
  BUF_X1 U967 ( .A(n1), .Z(n255) );
  BUF_X1 U968 ( .A(n46), .Z(n125) );
  BUF_X1 U969 ( .A(n45), .Z(n128) );
  BUF_X1 U970 ( .A(n44), .Z(n131) );
  BUF_X1 U971 ( .A(n43), .Z(n134) );
  BUF_X1 U972 ( .A(n42), .Z(n137) );
  BUF_X1 U973 ( .A(n41), .Z(n140) );
  BUF_X1 U974 ( .A(n15), .Z(n211) );
  BUF_X1 U975 ( .A(n16), .Z(n208) );
  BUF_X1 U976 ( .A(n14), .Z(n214) );
  BUF_X1 U977 ( .A(n13), .Z(n217) );
  BUF_X1 U978 ( .A(n12), .Z(n220) );
  BUF_X1 U979 ( .A(n11), .Z(n223) );
  BUF_X1 U980 ( .A(n10), .Z(n226) );
  BUF_X1 U981 ( .A(n9), .Z(n229) );
  BUF_X1 U982 ( .A(n8), .Z(n232) );
  BUF_X1 U983 ( .A(n7), .Z(n235) );
  BUF_X1 U984 ( .A(n21), .Z(n194) );
  BUF_X1 U985 ( .A(n22), .Z(n191) );
  BUF_X1 U986 ( .A(n20), .Z(n197) );
  BUF_X1 U987 ( .A(n19), .Z(n200) );
  BUF_X1 U988 ( .A(n14), .Z(n215) );
  BUF_X1 U989 ( .A(n13), .Z(n218) );
  BUF_X1 U990 ( .A(n18), .Z(n203) );
  BUF_X1 U991 ( .A(n17), .Z(n206) );
  BUF_X1 U992 ( .A(n16), .Z(n209) );
  BUF_X1 U993 ( .A(n15), .Z(n212) );
  BUF_X1 U994 ( .A(n12), .Z(n221) );
  BUF_X1 U995 ( .A(n11), .Z(n224) );
  BUF_X1 U996 ( .A(n10), .Z(n227) );
  BUF_X1 U997 ( .A(n9), .Z(n230) );
  BUF_X1 U998 ( .A(n8), .Z(n233) );
  BUF_X1 U999 ( .A(n7), .Z(n236) );
  BUF_X1 U1000 ( .A(n6), .Z(n239) );
  BUF_X1 U1001 ( .A(n5), .Z(n242) );
  BUF_X1 U1002 ( .A(n54), .Z(n100) );
  BUF_X2 U1003 ( .A(n28), .Z(n177) );
  BUF_X1 U1004 ( .A(n6), .Z(n238) );
  BUF_X1 U1005 ( .A(n4), .Z(n245) );
  BUF_X1 U1006 ( .A(n3), .Z(n248) );
  BUF_X1 U1007 ( .A(n48), .Z(n119) );
  BUF_X1 U1008 ( .A(n47), .Z(n122) );
  BUF_X1 U1009 ( .A(n44), .Z(n132) );
  BUF_X1 U1010 ( .A(n52), .Z(n108) );
  BUF_X1 U1011 ( .A(n50), .Z(n114) );
  BUF_X1 U1012 ( .A(n48), .Z(n120) );
  BUF_X1 U1013 ( .A(n43), .Z(n135) );
  BUF_X1 U1014 ( .A(n40), .Z(n144) );
  BUF_X1 U1015 ( .A(n38), .Z(n150) );
  BUF_X1 U1016 ( .A(n35), .Z(n159) );
  BUF_X1 U1017 ( .A(n53), .Z(n105) );
  BUF_X1 U1018 ( .A(n5), .Z(n241) );
  BUF_X2 U1019 ( .A(n31), .Z(n169) );
  BUF_X1 U1020 ( .A(n34), .Z(n162) );
  BUF_X2 U1021 ( .A(n30), .Z(n172) );
  BUF_X1 U1022 ( .A(shiftedA_62__63_), .Z(n342) );
  BUF_X2 U1023 ( .A(shiftedA_2__63_), .Z(n352) );
  BUF_X2 U1024 ( .A(shiftedA_5__63_), .Z(n361) );
  BUF_X2 U1025 ( .A(shiftedA_11__63_), .Z(n264) );
  BUF_X2 U1026 ( .A(shiftedA_63__63_), .Z(n343) );
  BUF_X2 U1027 ( .A(shiftedA_61__63_), .Z(n337) );
  BUF_X2 U1028 ( .A(shiftedA_62__63_), .Z(n340) );
  BUF_X2 U1029 ( .A(shiftedA_60__63_), .Z(n334) );
  BUF_X2 U1030 ( .A(shiftedA_59__63_), .Z(n331) );
  BUF_X2 U1031 ( .A(shiftedA_57__63_), .Z(n325) );
  BUF_X2 U1032 ( .A(shiftedA_54__63_), .Z(n316) );
  BUF_X2 U1033 ( .A(shiftedA_53__63_), .Z(n314) );
  BUF_X2 U1034 ( .A(shiftedA_0__63_), .Z(n347) );
  BUF_X2 U1035 ( .A(shiftedA_3__63_), .Z(n355) );
  BUF_X2 U1036 ( .A(shiftedA_6__63_), .Z(n364) );
  BUF_X2 U1037 ( .A(shiftedA_9__63_), .Z(n260) );
  BUF_X2 U1038 ( .A(shiftedA_12__63_), .Z(n266) );
  BUF_X2 U1039 ( .A(shiftedA_63__63_), .Z(n344) );
  BUF_X2 U1040 ( .A(shiftedA_62__63_), .Z(n341) );
  BUF_X2 U1041 ( .A(shiftedA_61__63_), .Z(n338) );
  BUF_X2 U1042 ( .A(shiftedA_60__63_), .Z(n335) );
  BUF_X2 U1043 ( .A(shiftedA_59__63_), .Z(n332) );
  BUF_X2 U1044 ( .A(shiftedA_57__63_), .Z(n326) );
  BUF_X2 U1045 ( .A(shiftedA_1__63_), .Z(n349) );
  BUF_X2 U1046 ( .A(shiftedA_4__63_), .Z(n358) );
  BUF_X2 U1047 ( .A(shiftedA_7__63_), .Z(n367) );
  BUF_X2 U1048 ( .A(shiftedA_10__63_), .Z(n262) );
  BUF_X1 U1049 ( .A(shiftedA_61__63_), .Z(n339) );
  BUF_X1 U1050 ( .A(shiftedA_60__63_), .Z(n336) );
  BUF_X1 U1051 ( .A(shiftedA_63__63_), .Z(n345) );
  BUF_X1 U1052 ( .A(shiftedA_51__63_), .Z(n311) );
  BUF_X1 U1053 ( .A(shiftedA_59__63_), .Z(n333) );
  BUF_X1 U1054 ( .A(n40), .Z(n143) );
  BUF_X1 U1055 ( .A(n39), .Z(n146) );
  BUF_X1 U1056 ( .A(n38), .Z(n149) );
  BUF_X1 U1057 ( .A(n37), .Z(n152) );
  BUF_X1 U1058 ( .A(n48), .Z(n118) );
  BUF_X1 U1059 ( .A(n35), .Z(n158) );
  BUF_X1 U1060 ( .A(n47), .Z(n121) );
  BUF_X1 U1061 ( .A(n36), .Z(n155) );
  BUF_X1 U1062 ( .A(n34), .Z(n161) );
  BUF_X1 U1063 ( .A(n46), .Z(n124) );
  BUF_X1 U1064 ( .A(n33), .Z(n164) );
  BUF_X1 U1065 ( .A(n45), .Z(n127) );
  BUF_X1 U1066 ( .A(n32), .Z(n167) );
  BUF_X1 U1067 ( .A(n44), .Z(n130) );
  BUF_X1 U1068 ( .A(n43), .Z(n133) );
  BUF_X1 U1069 ( .A(n42), .Z(n136) );
  BUF_X1 U1070 ( .A(n41), .Z(n139) );
  BUF_X1 U1071 ( .A(n40), .Z(n142) );
  BUF_X1 U1072 ( .A(n2), .Z(n251) );
  BUF_X1 U1073 ( .A(n1), .Z(n254) );
  BUF_X1 U1074 ( .A(n33), .Z(n165) );
  BUF_X1 U1075 ( .A(n32), .Z(n168) );
  BUF_X1 U1076 ( .A(n4), .Z(n244) );
  BUF_X1 U1077 ( .A(n3), .Z(n247) );
  BUF_X1 U1078 ( .A(n2), .Z(n250) );
  BUF_X1 U1079 ( .A(n1), .Z(n253) );
  BUF_X1 U1080 ( .A(shiftedA_57__63_), .Z(n327) );
  BUF_X1 U1081 ( .A(shiftedA_13__63_), .Z(n269) );
  BUF_X1 U1082 ( .A(shiftedA_1__63_), .Z(n351) );
  BUF_X1 U1083 ( .A(shiftedA_50__63_), .Z(n309) );
  BUF_X2 U1084 ( .A(shiftedA_2__63_), .Z(n353) );
  BUF_X2 U1085 ( .A(shiftedA_14__63_), .Z(n270) );
  BUF_X2 U1086 ( .A(shiftedA_5__63_), .Z(n362) );
  BUF_X2 U1087 ( .A(shiftedA_51__63_), .Z(n310) );
  BUF_X2 U1088 ( .A(shiftedA_52__63_), .Z(n312) );
  BUF_X2 U1089 ( .A(shiftedA_50__63_), .Z(n308) );
  BUF_X2 U1090 ( .A(shiftedA_49__63_), .Z(n306) );
  BUF_X2 U1091 ( .A(shiftedA_3__63_), .Z(n356) );
  BUF_X2 U1092 ( .A(shiftedA_6__63_), .Z(n365) );
  BUF_X2 U1093 ( .A(shiftedA_1__63_), .Z(n350) );
  BUF_X2 U1094 ( .A(shiftedA_4__63_), .Z(n359) );
  BUF_X2 U1095 ( .A(shiftedA_13__63_), .Z(n268) );
  BUF_X2 U1096 ( .A(shiftedA_7__63_), .Z(n368) );
  BUF_X1 U1097 ( .A(shiftedA_49__63_), .Z(n307) );
  BUF_X1 U1098 ( .A(shiftedA_0__63_), .Z(n348) );
  BUF_X1 U1099 ( .A(shiftedA_12__63_), .Z(n267) );
  BUF_X1 U1100 ( .A(n39), .Z(n145) );
  BUF_X1 U1101 ( .A(n38), .Z(n148) );
  BUF_X1 U1102 ( .A(n37), .Z(n151) );
  BUF_X1 U1103 ( .A(n35), .Z(n157) );
  BUF_X1 U1104 ( .A(n36), .Z(n154) );
  BUF_X1 U1105 ( .A(n34), .Z(n160) );
  BUF_X1 U1106 ( .A(n33), .Z(n163) );
  BUF_X1 U1107 ( .A(n32), .Z(n166) );
  BUF_X1 U1108 ( .A(shiftedA_14__63_), .Z(n271) );
  BUF_X1 U1109 ( .A(shiftedA_2__63_), .Z(n354) );
  BUF_X1 U1110 ( .A(shiftedA_3__63_), .Z(n357) );
  BUF_X1 U1111 ( .A(shiftedA_4__63_), .Z(n360) );
  BUF_X1 U1112 ( .A(shiftedA_5__63_), .Z(n363) );
  BUF_X1 U1113 ( .A(shiftedA_6__63_), .Z(n366) );
  AND2_X1 U1114 ( .A1(n372), .A2(n375), .ZN(shiftedA_32__63_) );
  BUF_X1 U1115 ( .A(shiftedA_7__63_), .Z(n369) );
  BUF_X1 U1116 ( .A(a[31]), .Z(n373) );
  INV_X1 U1117 ( .A(a[21]), .ZN(n10) );
  INV_X1 U1118 ( .A(a[22]), .ZN(n9) );
  INV_X1 U1119 ( .A(a[23]), .ZN(n8) );
  INV_X1 U1120 ( .A(a[24]), .ZN(n7) );
  INV_X1 U1121 ( .A(b[21]), .ZN(n41) );
  INV_X1 U1122 ( .A(b[23]), .ZN(n39) );
  INV_X1 U1123 ( .A(b[24]), .ZN(n38) );
  INV_X1 U1124 ( .A(a[9]), .ZN(n22) );
  INV_X1 U1125 ( .A(a[10]), .ZN(n21) );
  INV_X1 U1126 ( .A(b[9]), .ZN(n53) );
  INV_X1 U1127 ( .A(a[11]), .ZN(n20) );
  INV_X1 U1128 ( .A(a[12]), .ZN(n19) );
  INV_X1 U1129 ( .A(a[16]), .ZN(n15) );
  INV_X1 U1130 ( .A(a[15]), .ZN(n16) );
  INV_X1 U1131 ( .A(a[13]), .ZN(n18) );
  INV_X1 U1132 ( .A(a[18]), .ZN(n13) );
  INV_X1 U1133 ( .A(a[14]), .ZN(n17) );
  INV_X1 U1134 ( .A(a[17]), .ZN(n14) );
  INV_X1 U1135 ( .A(a[19]), .ZN(n12) );
  INV_X1 U1136 ( .A(a[27]), .ZN(n4) );
  INV_X1 U1137 ( .A(a[28]), .ZN(n3) );
  INV_X1 U1138 ( .A(a[26]), .ZN(n5) );
  INV_X1 U1139 ( .A(a[25]), .ZN(n6) );
  INV_X1 U1140 ( .A(a[29]), .ZN(n2) );
  INV_X1 U1141 ( .A(a[30]), .ZN(n1) );
  INV_X1 U1142 ( .A(a[20]), .ZN(n11) );
  INV_X1 U1143 ( .A(b[5]), .ZN(n57) );
  INV_X1 U1144 ( .A(b[6]), .ZN(n56) );
  INV_X1 U1145 ( .A(b[7]), .ZN(n55) );
  INV_X1 U1146 ( .A(b[8]), .ZN(n54) );
  INV_X1 U1147 ( .A(b[12]), .ZN(n50) );
  INV_X1 U1148 ( .A(b[11]), .ZN(n51) );
  INV_X1 U1149 ( .A(b[10]), .ZN(n52) );
  INV_X1 U1150 ( .A(b[18]), .ZN(n44) );
  INV_X1 U1151 ( .A(b[13]), .ZN(n49) );
  INV_X1 U1152 ( .A(b[17]), .ZN(n45) );
  INV_X1 U1153 ( .A(b[14]), .ZN(n48) );
  INV_X1 U1154 ( .A(b[15]), .ZN(n47) );
  INV_X1 U1155 ( .A(b[16]), .ZN(n46) );
  INV_X1 U1156 ( .A(b[19]), .ZN(n43) );
  INV_X1 U1157 ( .A(b[20]), .ZN(n42) );
  INV_X1 U1158 ( .A(b[22]), .ZN(n40) );
  INV_X1 U1159 ( .A(b[25]), .ZN(n37) );
  INV_X1 U1160 ( .A(b[27]), .ZN(n35) );
  INV_X1 U1161 ( .A(b[26]), .ZN(n36) );
  INV_X1 U1162 ( .A(b[28]), .ZN(n34) );
  INV_X1 U1163 ( .A(b[2]), .ZN(n60) );
  BUF_X1 U1164 ( .A(a[31]), .Z(n374) );
  BUF_X1 U1165 ( .A(b[31]), .Z(n371) );
  BUF_X1 U1166 ( .A(b[31]), .Z(n370) );
  BUF_X1 U1167 ( .A(a[31]), .Z(n375) );
  AND2_X1 U1168 ( .A1(b[2]), .A2(n374), .ZN(shiftedA_2__63_) );
  AND2_X1 U1169 ( .A1(n370), .A2(a[3]), .ZN(shiftedA_60__63_) );
  AND2_X1 U1170 ( .A1(b[5]), .A2(n375), .ZN(shiftedA_5__63_) );
  AND2_X1 U1171 ( .A1(b[6]), .A2(n375), .ZN(shiftedA_6__63_) );
  AND2_X1 U1172 ( .A1(b[7]), .A2(n375), .ZN(shiftedA_7__63_) );
  INV_X1 U1173 ( .A(b[29]), .ZN(n33) );
  INV_X1 U1174 ( .A(b[30]), .ZN(n32) );
  AND2_X1 U1175 ( .A1(n371), .A2(a[12]), .ZN(shiftedA_51__63_) );
  AND2_X1 U1176 ( .A1(b[10]), .A2(n373), .ZN(shiftedA_10__63_) );
  AND2_X1 U1177 ( .A1(b[11]), .A2(n373), .ZN(shiftedA_11__63_) );
  AND2_X1 U1178 ( .A1(b[12]), .A2(n373), .ZN(shiftedA_12__63_) );
  AND2_X1 U1179 ( .A1(n370), .A2(a[9]), .ZN(shiftedA_54__63_) );
  AND2_X1 U1180 ( .A1(n370), .A2(a[10]), .ZN(shiftedA_53__63_) );
  AND2_X1 U1181 ( .A1(n370), .A2(a[11]), .ZN(shiftedA_52__63_) );
  AND2_X1 U1182 ( .A1(n375), .A2(b[9]), .ZN(shiftedA_9__63_) );
  AND2_X1 U1183 ( .A1(b[8]), .A2(n375), .ZN(shiftedA_8__63_) );
  AND2_X1 U1184 ( .A1(n370), .A2(a[8]), .ZN(shiftedA_55__63_) );
  AND2_X1 U1185 ( .A1(n372), .A2(a[24]), .ZN(shiftedA_39__63_) );
  BUF_X1 U1186 ( .A(b[31]), .Z(n372) );
  AND2_X1 U1187 ( .A1(n371), .A2(a[13]), .ZN(shiftedA_50__63_) );
  AND2_X1 U1188 ( .A1(n371), .A2(a[14]), .ZN(shiftedA_49__63_) );
  AND2_X1 U1189 ( .A1(b[13]), .A2(n373), .ZN(shiftedA_13__63_) );
  AND2_X1 U1190 ( .A1(b[14]), .A2(n373), .ZN(shiftedA_14__63_) );
  AND2_X1 U1191 ( .A1(n371), .A2(a[19]), .ZN(shiftedA_44__63_) );
  AND2_X1 U1192 ( .A1(n371), .A2(a[15]), .ZN(shiftedA_48__63_) );
  AND2_X1 U1193 ( .A1(n371), .A2(a[16]), .ZN(shiftedA_47__63_) );
  AND2_X1 U1194 ( .A1(n371), .A2(a[18]), .ZN(shiftedA_45__63_) );
  AND2_X1 U1195 ( .A1(n371), .A2(a[20]), .ZN(shiftedA_43__63_) );
  AND2_X1 U1196 ( .A1(n371), .A2(a[17]), .ZN(shiftedA_46__63_) );
  AND2_X1 U1197 ( .A1(b[20]), .A2(n374), .ZN(shiftedA_20__63_) );
  AND2_X1 U1198 ( .A1(b[15]), .A2(n373), .ZN(shiftedA_15__63_) );
  AND2_X1 U1199 ( .A1(b[16]), .A2(n373), .ZN(shiftedA_16__63_) );
  AND2_X1 U1200 ( .A1(b[17]), .A2(n373), .ZN(shiftedA_17__63_) );
  AND2_X1 U1201 ( .A1(b[18]), .A2(n373), .ZN(shiftedA_18__63_) );
  AND2_X1 U1202 ( .A1(b[19]), .A2(n373), .ZN(shiftedA_19__63_) );
  AND2_X1 U1203 ( .A1(n372), .A2(a[25]), .ZN(shiftedA_38__63_) );
  AND2_X1 U1204 ( .A1(b[25]), .A2(n374), .ZN(shiftedA_25__63_) );
  AND2_X1 U1205 ( .A1(b[26]), .A2(n374), .ZN(shiftedA_26__63_) );
  AND2_X1 U1206 ( .A1(n372), .A2(a[26]), .ZN(shiftedA_37__63_) );
  AND2_X1 U1207 ( .A1(b[27]), .A2(n374), .ZN(shiftedA_27__63_) );
  AND2_X1 U1208 ( .A1(n372), .A2(a[27]), .ZN(shiftedA_36__63_) );
  AND2_X1 U1209 ( .A1(n372), .A2(a[28]), .ZN(shiftedA_35__63_) );
  AND2_X1 U1210 ( .A1(b[28]), .A2(n374), .ZN(shiftedA_28__63_) );
  AND2_X1 U1211 ( .A1(b[24]), .A2(n374), .ZN(shiftedA_24__63_) );
  AND2_X1 U1212 ( .A1(b[29]), .A2(n374), .ZN(shiftedA_29__63_) );
  AND2_X1 U1213 ( .A1(n372), .A2(a[29]), .ZN(shiftedA_34__63_) );
  AND2_X1 U1214 ( .A1(b[30]), .A2(n374), .ZN(shiftedA_30__63_) );
  AND2_X1 U1215 ( .A1(n372), .A2(a[30]), .ZN(shiftedA_33__63_) );
  INV_X1 U1216 ( .A(a[0]), .ZN(n31) );
  AND2_X1 U1217 ( .A1(n370), .A2(a[0]), .ZN(shiftedA_63__63_) );
  CLKBUF_X1 U1219 ( .A(n68), .Z(n89) );
  NOR2_X1 U1220 ( .A1(n181), .A2(n165), .ZN(shiftedA_29__34_) );
  NOR2_X1 U1221 ( .A1(n181), .A2(n168), .ZN(shiftedA_30__35_) );
  NOR2_X1 U1222 ( .A1(n181), .A2(n162), .ZN(shiftedA_28__33_) );
  NOR2_X1 U1223 ( .A1(n181), .A2(n159), .ZN(shiftedA_27__32_) );
  NOR2_X1 U1224 ( .A1(n181), .A2(n102), .ZN(shiftedA_8__13_) );
  NOR2_X1 U1225 ( .A1(n105), .A2(n181), .ZN(shiftedA_9__14_) );
  NOR2_X1 U1226 ( .A1(n181), .A2(n99), .ZN(shiftedA_7__12_) );
  NOR2_X1 U1227 ( .A1(n181), .A2(n93), .ZN(shiftedA_5__10_) );
  NOR2_X1 U1228 ( .A1(n181), .A2(n96), .ZN(shiftedA_6__11_) );
  NOR2_X1 U1229 ( .A1(n73), .A2(n84), .ZN(shiftedA_2__7_) );
  NOR2_X1 U1230 ( .A1(n188), .A2(n122), .ZN(shiftedA_15__23_) );
  NOR2_X1 U1231 ( .A1(n187), .A2(n119), .ZN(shiftedA_14__22_) );
  NOR2_X1 U1232 ( .A1(n188), .A2(n116), .ZN(shiftedA_13__21_) );
  NOR2_X1 U1233 ( .A1(n187), .A2(n110), .ZN(shiftedA_11__19_) );
  NOR2_X1 U1234 ( .A1(n188), .A2(n113), .ZN(shiftedA_12__20_) );
  NOR2_X1 U1235 ( .A1(n187), .A2(n107), .ZN(shiftedA_10__18_) );
  CLKBUF_X1 U1236 ( .A(n24), .Z(n186) );
  INV_X1 U1237 ( .A(b[3]), .ZN(n75) );
  NOR2_X1 U1238 ( .A1(n181), .A2(n156), .ZN(shiftedA_26__31_) );
  NOR2_X1 U1239 ( .A1(n181), .A2(n153), .ZN(shiftedA_25__30_) );
  NOR2_X1 U1240 ( .A1(n181), .A2(n150), .ZN(shiftedA_24__29_) );
  NOR2_X1 U1241 ( .A1(n181), .A2(n147), .ZN(shiftedA_23__28_) );
  NOR2_X1 U1242 ( .A1(n181), .A2(n144), .ZN(shiftedA_22__27_) );
  NOR2_X1 U1243 ( .A1(n181), .A2(n138), .ZN(shiftedA_20__25_) );
  NOR2_X1 U1244 ( .A1(n181), .A2(n141), .ZN(shiftedA_21__26_) );
  NOR2_X1 U1245 ( .A1(n181), .A2(n135), .ZN(shiftedA_19__24_) );
  NOR2_X1 U1246 ( .A1(n181), .A2(n129), .ZN(shiftedA_17__22_) );
  NOR2_X1 U1247 ( .A1(n181), .A2(n132), .ZN(shiftedA_18__23_) );
  NOR2_X1 U1248 ( .A1(n181), .A2(n126), .ZN(shiftedA_16__21_) );
  AND2_X1 U1249 ( .A1(n370), .A2(n66), .ZN(shiftedA_59__63_) );
  NOR2_X1 U1250 ( .A1(n79), .A2(n162), .ZN(shiftedA_28__31_) );
  NOR2_X1 U1251 ( .A1(n79), .A2(n150), .ZN(shiftedA_24__27_) );
  NOR2_X1 U1252 ( .A1(n79), .A2(n144), .ZN(shiftedA_22__25_) );
  NOR2_X1 U1253 ( .A1(n79), .A2(n135), .ZN(shiftedA_19__22_) );
  NOR2_X1 U1254 ( .A1(n79), .A2(n132), .ZN(shiftedA_18__21_) );
  NOR2_X1 U1255 ( .A1(n79), .A2(n120), .ZN(shiftedA_14__17_) );
  NOR2_X1 U1256 ( .A1(n79), .A2(n114), .ZN(shiftedA_12__15_) );
  NOR2_X1 U1257 ( .A1(n79), .A2(n108), .ZN(shiftedA_10__13_) );
  NOR2_X1 U1258 ( .A1(n79), .A2(n84), .ZN(shiftedA_2__5_) );
  CLKBUF_X1 U1259 ( .A(n183), .Z(n78) );
  INV_X1 U1260 ( .A(a[8]), .ZN(n23) );
  AND2_X1 U1261 ( .A1(n370), .A2(a[5]), .ZN(shiftedA_58__63_) );
  NOR2_X1 U1262 ( .A1(n179), .A2(n162), .ZN(shiftedA_28__32_) );
  NOR2_X1 U1263 ( .A1(n179), .A2(n150), .ZN(shiftedA_24__28_) );
  NOR2_X1 U1264 ( .A1(n180), .A2(n144), .ZN(shiftedA_22__26_) );
  NOR2_X1 U1265 ( .A1(n180), .A2(n135), .ZN(shiftedA_19__23_) );
  NOR2_X1 U1266 ( .A1(n180), .A2(n132), .ZN(shiftedA_18__22_) );
  NOR2_X1 U1267 ( .A1(n180), .A2(n120), .ZN(shiftedA_14__18_) );
  NOR2_X1 U1268 ( .A1(n180), .A2(n114), .ZN(shiftedA_12__16_) );
  NOR2_X1 U1269 ( .A1(n180), .A2(n108), .ZN(shiftedA_10__14_) );
  NOR2_X1 U1270 ( .A1(n180), .A2(n84), .ZN(shiftedA_2__6_) );
  NOR2_X1 U1271 ( .A1(n192), .A2(n67), .ZN(shiftedA_0__9_) );
  NOR2_X1 U1272 ( .A1(n189), .A2(n67), .ZN(shiftedA_0__8_) );
  NOR2_X1 U1273 ( .A1(n62), .A2(n25), .ZN(shiftedA_0__6_) );
  NOR2_X1 U1274 ( .A1(n179), .A2(n67), .ZN(shiftedA_0__4_) );
  NOR2_X1 U1275 ( .A1(n79), .A2(n80), .ZN(shiftedA_0__3_) );
  NOR2_X1 U1276 ( .A1(n255), .A2(n67), .ZN(shiftedA_0__30_) );
  NOR2_X1 U1277 ( .A1(n176), .A2(n80), .ZN(shiftedA_0__2_) );
  NOR2_X1 U1278 ( .A1(n252), .A2(n80), .ZN(shiftedA_0__29_) );
  NOR2_X1 U1279 ( .A1(n249), .A2(n80), .ZN(shiftedA_0__28_) );
  NOR2_X1 U1280 ( .A1(n246), .A2(n80), .ZN(shiftedA_0__27_) );
  AND2_X1 U1281 ( .A1(n66), .A2(b[3]), .ZN(shiftedA_3__7_) );
  INV_X1 U1282 ( .A(a[1]), .ZN(n30) );
  AND2_X1 U1283 ( .A1(n370), .A2(a[1]), .ZN(shiftedA_62__63_) );
  AND2_X1 U1284 ( .A1(a[3]), .A2(b[4]), .ZN(shiftedA_4__7_) );
  NOR2_X1 U1285 ( .A1(n76), .A2(n168), .ZN(shiftedA_30__32_) );
  NOR2_X1 U1286 ( .A1(n76), .A2(n165), .ZN(shiftedA_29__31_) );
  AND2_X1 U1287 ( .A1(n370), .A2(a[2]), .ZN(shiftedA_61__63_) );
  NOR2_X1 U1288 ( .A1(n76), .A2(n162), .ZN(shiftedA_28__30_) );
  NOR2_X1 U1289 ( .A1(n76), .A2(n159), .ZN(shiftedA_27__29_) );
  NOR2_X1 U1290 ( .A1(n176), .A2(n102), .ZN(shiftedA_8__10_) );
  NOR2_X1 U1291 ( .A1(n63), .A2(n97), .ZN(shiftedA_7__9_) );
  NOR2_X1 U1292 ( .A1(n63), .A2(n84), .ZN(shiftedA_2__4_) );
  NOR2_X1 U1293 ( .A1(n105), .A2(n63), .ZN(shiftedA_9__11_) );
  NOR2_X1 U1294 ( .A1(n29), .A2(n91), .ZN(shiftedA_5__7_) );
  NOR2_X1 U1295 ( .A1(n172), .A2(n165), .ZN(shiftedA_29__30_) );
  NOR2_X1 U1296 ( .A1(n172), .A2(n168), .ZN(shiftedA_30__31_) );
  NOR2_X1 U1297 ( .A1(n172), .A2(n162), .ZN(shiftedA_28__29_) );
  NOR2_X1 U1298 ( .A1(n172), .A2(n159), .ZN(shiftedA_27__28_) );
  NOR2_X1 U1299 ( .A1(n172), .A2(n100), .ZN(shiftedA_8__9_) );
  NOR2_X1 U1300 ( .A1(n172), .A2(n84), .ZN(shiftedA_2__3_) );
  NOR2_X1 U1301 ( .A1(n172), .A2(n97), .ZN(shiftedA_7__8_) );
  NOR2_X1 U1302 ( .A1(n172), .A2(n91), .ZN(shiftedA_5__6_) );
  NOR2_X1 U1303 ( .A1(n172), .A2(n94), .ZN(shiftedA_6__7_) );
  NOR2_X1 U1304 ( .A1(n105), .A2(n172), .ZN(shiftedA_9__10_) );
  NOR2_X1 U1305 ( .A1(n181), .A2(n123), .ZN(shiftedA_15__20_) );
  NOR2_X1 U1306 ( .A1(n181), .A2(n120), .ZN(shiftedA_14__19_) );
  NOR2_X1 U1307 ( .A1(n181), .A2(n117), .ZN(shiftedA_13__18_) );
  NOR2_X1 U1308 ( .A1(n181), .A2(n111), .ZN(shiftedA_11__16_) );
  NOR2_X1 U1309 ( .A1(n181), .A2(n114), .ZN(shiftedA_12__17_) );
  NOR2_X1 U1310 ( .A1(n181), .A2(n108), .ZN(shiftedA_10__15_) );
  INV_X1 U1311 ( .A(a[4]), .ZN(n27) );
  BUF_X2 U1312 ( .A(n28), .Z(n79) );
  INV_X1 U1313 ( .A(a[3]), .ZN(n28) );
  AND2_X1 U1314 ( .A1(n370), .A2(a[6]), .ZN(shiftedA_57__63_) );
  INV_X1 U1315 ( .A(a[6]), .ZN(n25) );
  AND2_X1 U1316 ( .A1(n370), .A2(a[7]), .ZN(shiftedA_56__63_) );
  NOR2_X1 U1317 ( .A1(n185), .A2(n122), .ZN(shiftedA_15__22_) );
  NOR2_X1 U1318 ( .A1(n184), .A2(n119), .ZN(shiftedA_14__21_) );
  NOR2_X1 U1319 ( .A1(n77), .A2(n116), .ZN(shiftedA_13__20_) );
  NOR2_X1 U1320 ( .A1(n185), .A2(n110), .ZN(shiftedA_11__18_) );
  NOR2_X1 U1321 ( .A1(n184), .A2(n113), .ZN(shiftedA_12__19_) );
  NOR2_X1 U1322 ( .A1(n184), .A2(n107), .ZN(shiftedA_10__17_) );
  INV_X1 U1323 ( .A(a[7]), .ZN(n24) );
  AND2_X1 U1324 ( .A1(n71), .A2(n373), .ZN(shiftedA_0__63_) );
  NOR2_X1 U1325 ( .A1(n254), .A2(n82), .ZN(shiftedA_1__31_) );
  AND2_X1 U1326 ( .A1(n64), .A2(n373), .ZN(shiftedA_1__63_) );
  NOR2_X1 U1327 ( .A1(n251), .A2(n82), .ZN(shiftedA_1__30_) );
  NOR2_X1 U1328 ( .A1(n248), .A2(n82), .ZN(shiftedA_1__29_) );
  NOR2_X1 U1329 ( .A1(n245), .A2(n82), .ZN(shiftedA_1__28_) );
  NOR2_X1 U1330 ( .A1(n173), .A2(n82), .ZN(shiftedA_1__2_) );
  NOR2_X1 U1331 ( .A1(n63), .A2(n82), .ZN(shiftedA_1__3_) );
  NOR2_X1 U1332 ( .A1(n189), .A2(n61), .ZN(shiftedA_1__9_) );
  NOR2_X1 U1333 ( .A1(n79), .A2(n61), .ZN(shiftedA_1__4_) );
  NOR2_X1 U1334 ( .A1(n186), .A2(n61), .ZN(shiftedA_1__8_) );
  NOR2_X1 U1335 ( .A1(n253), .A2(n88), .ZN(shiftedA_3__33_) );
  AND2_X1 U1336 ( .A1(n69), .A2(n375), .ZN(shiftedA_3__63_) );
  NOR2_X1 U1337 ( .A1(n250), .A2(n87), .ZN(shiftedA_3__32_) );
  NOR2_X1 U1338 ( .A1(n247), .A2(n88), .ZN(shiftedA_3__31_) );
  NOR2_X1 U1339 ( .A1(n244), .A2(n87), .ZN(shiftedA_3__30_) );
  NOR2_X1 U1340 ( .A1(n241), .A2(n88), .ZN(shiftedA_3__29_) );
  NOR2_X1 U1341 ( .A1(n169), .A2(n87), .ZN(shiftedA_3__3_) );
  NOR2_X1 U1342 ( .A1(n172), .A2(n87), .ZN(shiftedA_3__4_) );
  NOR2_X1 U1343 ( .A1(n25), .A2(n75), .ZN(shiftedA_3__9_) );
  NOR2_X1 U1344 ( .A1(n28), .A2(n75), .ZN(shiftedA_3__6_) );
  NOR2_X1 U1345 ( .A1(n72), .A2(n75), .ZN(shiftedA_3__5_) );
  NOR2_X1 U1346 ( .A1(n73), .A2(n75), .ZN(shiftedA_3__8_) );
  INV_X1 U1347 ( .A(b[3]), .ZN(n59) );
  NOR2_X1 U1348 ( .A1(n253), .A2(n58), .ZN(shiftedA_4__34_) );
  AND2_X1 U1349 ( .A1(n70), .A2(n375), .ZN(shiftedA_4__63_) );
  NOR2_X1 U1350 ( .A1(n250), .A2(n90), .ZN(shiftedA_4__33_) );
  NOR2_X1 U1351 ( .A1(n247), .A2(n90), .ZN(shiftedA_4__32_) );
  NOR2_X1 U1352 ( .A1(n244), .A2(n90), .ZN(shiftedA_4__31_) );
  NOR2_X1 U1353 ( .A1(n241), .A2(n90), .ZN(shiftedA_4__30_) );
  NOR2_X1 U1354 ( .A1(n238), .A2(n90), .ZN(shiftedA_4__29_) );
  NOR2_X1 U1355 ( .A1(n169), .A2(n58), .ZN(shiftedA_4__4_) );
  NOR2_X1 U1356 ( .A1(n73), .A2(n58), .ZN(shiftedA_4__9_) );
  NOR2_X1 U1357 ( .A1(n30), .A2(n58), .ZN(shiftedA_4__5_) );
  NOR2_X1 U1358 ( .A1(n73), .A2(n67), .ZN(shiftedA_0__5_) );
  NOR2_X1 U1359 ( .A1(n27), .A2(n61), .ZN(shiftedA_1__5_) );
  BUF_X1 U1360 ( .A(shiftedA_8__63_), .Z(n256) );
  BUF_X1 U1361 ( .A(shiftedA_8__63_), .Z(n257) );
  BUF_X1 U1362 ( .A(shiftedA_8__63_), .Z(n258) );
  BUF_X1 U1363 ( .A(shiftedA_8__63_), .Z(n259) );
  BUF_X1 U1364 ( .A(shiftedA_15__63_), .Z(n272) );
  BUF_X1 U1365 ( .A(shiftedA_15__63_), .Z(n273) );
  BUF_X1 U1366 ( .A(shiftedA_15__63_), .Z(n274) );
  BUF_X1 U1367 ( .A(shiftedA_16__63_), .Z(n275) );
  BUF_X1 U1368 ( .A(shiftedA_16__63_), .Z(n276) );
  BUF_X1 U1369 ( .A(shiftedA_16__63_), .Z(n277) );
  BUF_X1 U1370 ( .A(shiftedA_17__63_), .Z(n278) );
  BUF_X1 U1371 ( .A(shiftedA_17__63_), .Z(n279) );
  BUF_X1 U1372 ( .A(shiftedA_17__63_), .Z(n280) );
  BUF_X1 U1373 ( .A(shiftedA_18__63_), .Z(n281) );
  BUF_X1 U1374 ( .A(shiftedA_18__63_), .Z(n282) );
  BUF_X1 U1375 ( .A(shiftedA_18__63_), .Z(n283) );
  BUF_X1 U1376 ( .A(shiftedA_19__63_), .Z(n284) );
  BUF_X1 U1377 ( .A(shiftedA_19__63_), .Z(n285) );
  BUF_X1 U1378 ( .A(shiftedA_19__63_), .Z(n286) );
  BUF_X1 U1379 ( .A(shiftedA_20__63_), .Z(n287) );
  BUF_X1 U1380 ( .A(shiftedA_20__63_), .Z(n288) );
  BUF_X1 U1381 ( .A(shiftedA_43__63_), .Z(n289) );
  BUF_X1 U1382 ( .A(shiftedA_43__63_), .Z(n290) );
  BUF_X1 U1383 ( .A(shiftedA_44__63_), .Z(n291) );
  BUF_X1 U1384 ( .A(shiftedA_44__63_), .Z(n292) );
  BUF_X1 U1385 ( .A(shiftedA_44__63_), .Z(n293) );
  BUF_X1 U1386 ( .A(shiftedA_45__63_), .Z(n294) );
  BUF_X1 U1387 ( .A(shiftedA_45__63_), .Z(n295) );
  BUF_X1 U1388 ( .A(shiftedA_45__63_), .Z(n296) );
  BUF_X1 U1389 ( .A(shiftedA_46__63_), .Z(n297) );
  BUF_X1 U1390 ( .A(shiftedA_46__63_), .Z(n298) );
  BUF_X1 U1391 ( .A(shiftedA_46__63_), .Z(n299) );
  BUF_X1 U1392 ( .A(shiftedA_47__63_), .Z(n300) );
  BUF_X1 U1393 ( .A(shiftedA_47__63_), .Z(n301) );
  BUF_X1 U1394 ( .A(shiftedA_47__63_), .Z(n302) );
  BUF_X1 U1395 ( .A(shiftedA_48__63_), .Z(n303) );
  BUF_X1 U1396 ( .A(shiftedA_48__63_), .Z(n304) );
  BUF_X1 U1397 ( .A(shiftedA_48__63_), .Z(n305) );
  BUF_X1 U1398 ( .A(shiftedA_55__63_), .Z(n318) );
  BUF_X1 U1399 ( .A(shiftedA_55__63_), .Z(n319) );
  BUF_X1 U1400 ( .A(shiftedA_55__63_), .Z(n320) );
  BUF_X1 U1401 ( .A(shiftedA_55__63_), .Z(n321) );
endmodule


module regN_N64 ( clk, reset, in, out );
  input [63:0] in;
  output [63:0] out;
  input clk, reset;
  wire   n65, n64;

  DFF_X1 out_reg_63_ ( .D(n64), .CK(clk), .Q(out[63]) );
  SDFF_X1 out_reg_7_ ( .D(1'b0), .SI(n65), .SE(in[7]), .CK(clk), .Q(out[7]) );
  SDFF_X1 out_reg_8_ ( .D(1'b0), .SI(n65), .SE(in[8]), .CK(clk), .Q(out[8]) );
  SDFF_X1 out_reg_6_ ( .D(1'b0), .SI(n65), .SE(in[6]), .CK(clk), .Q(out[6]) );
  SDFF_X1 out_reg_9_ ( .D(1'b0), .SI(n65), .SE(in[9]), .CK(clk), .Q(out[9]) );
  SDFF_X1 out_reg_5_ ( .D(1'b0), .SI(n65), .SE(in[5]), .CK(clk), .Q(out[5]) );
  SDFF_X1 out_reg_10_ ( .D(1'b0), .SI(n65), .SE(in[10]), .CK(clk), .Q(out[10])
         );
  SDFF_X1 out_reg_11_ ( .D(1'b0), .SI(n65), .SE(in[11]), .CK(clk), .Q(out[11])
         );
  SDFF_X1 out_reg_0_ ( .D(1'b0), .SI(n65), .SE(in[0]), .CK(clk), .Q(out[0]) );
  SDFF_X1 out_reg_4_ ( .D(1'b0), .SI(n65), .SE(in[4]), .CK(clk), .Q(out[4]) );
  SDFF_X1 out_reg_3_ ( .D(1'b0), .SI(n65), .SE(in[3]), .CK(clk), .Q(out[3]) );
  SDFF_X1 out_reg_1_ ( .D(1'b0), .SI(n65), .SE(in[1]), .CK(clk), .Q(out[1]) );
  SDFF_X1 out_reg_12_ ( .D(1'b0), .SI(n65), .SE(in[12]), .CK(clk), .Q(out[12])
         );
  SDFF_X1 out_reg_2_ ( .D(1'b0), .SI(n65), .SE(in[2]), .CK(clk), .Q(out[2]) );
  SDFF_X1 out_reg_13_ ( .D(1'b0), .SI(n65), .SE(in[13]), .CK(clk), .Q(out[13])
         );
  SDFF_X1 out_reg_14_ ( .D(1'b0), .SI(n65), .SE(in[14]), .CK(clk), .Q(out[14])
         );
  SDFF_X1 out_reg_15_ ( .D(1'b0), .SI(n65), .SE(in[15]), .CK(clk), .Q(out[15])
         );
  SDFF_X1 out_reg_16_ ( .D(1'b0), .SI(n65), .SE(in[16]), .CK(clk), .Q(out[16])
         );
  SDFF_X1 out_reg_17_ ( .D(1'b0), .SI(n65), .SE(in[17]), .CK(clk), .Q(out[17])
         );
  SDFF_X1 out_reg_18_ ( .D(1'b0), .SI(n65), .SE(in[18]), .CK(clk), .Q(out[18])
         );
  SDFF_X1 out_reg_19_ ( .D(1'b0), .SI(n65), .SE(in[19]), .CK(clk), .Q(out[19])
         );
  SDFF_X1 out_reg_20_ ( .D(1'b0), .SI(n65), .SE(in[20]), .CK(clk), .Q(out[20])
         );
  SDFF_X1 out_reg_21_ ( .D(1'b0), .SI(n65), .SE(in[21]), .CK(clk), .Q(out[21])
         );
  SDFF_X1 out_reg_22_ ( .D(1'b0), .SI(n65), .SE(in[22]), .CK(clk), .Q(out[22])
         );
  SDFF_X1 out_reg_23_ ( .D(1'b0), .SI(n65), .SE(in[23]), .CK(clk), .Q(out[23])
         );
  SDFF_X1 out_reg_24_ ( .D(1'b0), .SI(n65), .SE(in[24]), .CK(clk), .Q(out[24])
         );
  SDFF_X1 out_reg_25_ ( .D(1'b0), .SI(n65), .SE(in[25]), .CK(clk), .Q(out[25])
         );
  SDFF_X1 out_reg_26_ ( .D(1'b0), .SI(n65), .SE(in[26]), .CK(clk), .Q(out[26])
         );
  SDFF_X1 out_reg_27_ ( .D(1'b0), .SI(n65), .SE(in[27]), .CK(clk), .Q(out[27])
         );
  SDFF_X1 out_reg_28_ ( .D(1'b0), .SI(n65), .SE(in[28]), .CK(clk), .Q(out[28])
         );
  SDFF_X1 out_reg_29_ ( .D(1'b0), .SI(n65), .SE(in[29]), .CK(clk), .Q(out[29])
         );
  SDFF_X1 out_reg_30_ ( .D(1'b0), .SI(n65), .SE(in[30]), .CK(clk), .Q(out[30])
         );
  SDFF_X1 out_reg_31_ ( .D(1'b0), .SI(n65), .SE(in[31]), .CK(clk), .Q(out[31])
         );
  SDFF_X1 out_reg_32_ ( .D(1'b0), .SI(n65), .SE(in[32]), .CK(clk), .Q(out[32])
         );
  SDFF_X1 out_reg_33_ ( .D(1'b0), .SI(n65), .SE(in[33]), .CK(clk), .Q(out[33])
         );
  SDFF_X1 out_reg_34_ ( .D(1'b0), .SI(n65), .SE(in[34]), .CK(clk), .Q(out[34])
         );
  SDFF_X1 out_reg_35_ ( .D(1'b0), .SI(n65), .SE(in[35]), .CK(clk), .Q(out[35])
         );
  SDFF_X1 out_reg_36_ ( .D(1'b0), .SI(n65), .SE(in[36]), .CK(clk), .Q(out[36])
         );
  SDFF_X1 out_reg_37_ ( .D(1'b0), .SI(n65), .SE(in[37]), .CK(clk), .Q(out[37])
         );
  SDFF_X1 out_reg_38_ ( .D(1'b0), .SI(n65), .SE(in[38]), .CK(clk), .Q(out[38])
         );
  SDFF_X1 out_reg_39_ ( .D(1'b0), .SI(n65), .SE(in[39]), .CK(clk), .Q(out[39])
         );
  SDFF_X1 out_reg_40_ ( .D(1'b0), .SI(n65), .SE(in[40]), .CK(clk), .Q(out[40])
         );
  SDFF_X1 out_reg_41_ ( .D(1'b0), .SI(n65), .SE(in[41]), .CK(clk), .Q(out[41])
         );
  SDFF_X1 out_reg_42_ ( .D(1'b0), .SI(n65), .SE(in[42]), .CK(clk), .Q(out[42])
         );
  SDFF_X1 out_reg_43_ ( .D(1'b0), .SI(n65), .SE(in[43]), .CK(clk), .Q(out[43])
         );
  SDFF_X1 out_reg_44_ ( .D(1'b0), .SI(n65), .SE(in[44]), .CK(clk), .Q(out[44])
         );
  SDFF_X1 out_reg_45_ ( .D(1'b0), .SI(n65), .SE(in[45]), .CK(clk), .Q(out[45])
         );
  SDFF_X1 out_reg_46_ ( .D(1'b0), .SI(n65), .SE(in[46]), .CK(clk), .Q(out[46])
         );
  SDFF_X1 out_reg_47_ ( .D(1'b0), .SI(n65), .SE(in[47]), .CK(clk), .Q(out[47])
         );
  SDFF_X1 out_reg_48_ ( .D(1'b0), .SI(n65), .SE(in[48]), .CK(clk), .Q(out[48])
         );
  SDFF_X1 out_reg_49_ ( .D(1'b0), .SI(n65), .SE(in[49]), .CK(clk), .Q(out[49])
         );
  SDFF_X1 out_reg_50_ ( .D(1'b0), .SI(n65), .SE(in[50]), .CK(clk), .Q(out[50])
         );
  SDFF_X1 out_reg_51_ ( .D(1'b0), .SI(n65), .SE(in[51]), .CK(clk), .Q(out[51])
         );
  SDFF_X1 out_reg_52_ ( .D(1'b0), .SI(n65), .SE(in[52]), .CK(clk), .Q(out[52])
         );
  SDFF_X1 out_reg_53_ ( .D(1'b0), .SI(n65), .SE(in[53]), .CK(clk), .Q(out[53])
         );
  SDFF_X1 out_reg_54_ ( .D(1'b0), .SI(n65), .SE(in[54]), .CK(clk), .Q(out[54])
         );
  SDFF_X1 out_reg_55_ ( .D(1'b0), .SI(n65), .SE(in[55]), .CK(clk), .Q(out[55])
         );
  SDFF_X1 out_reg_56_ ( .D(1'b0), .SI(n65), .SE(in[56]), .CK(clk), .Q(out[56])
         );
  SDFF_X1 out_reg_57_ ( .D(1'b0), .SI(n65), .SE(in[57]), .CK(clk), .Q(out[57])
         );
  SDFF_X1 out_reg_58_ ( .D(1'b0), .SI(n65), .SE(in[58]), .CK(clk), .Q(out[58])
         );
  SDFF_X1 out_reg_59_ ( .D(1'b0), .SI(n65), .SE(in[59]), .CK(clk), .Q(out[59])
         );
  SDFF_X1 out_reg_60_ ( .D(1'b0), .SI(n65), .SE(in[60]), .CK(clk), .Q(out[60])
         );
  SDFF_X1 out_reg_61_ ( .D(1'b0), .SI(n65), .SE(in[61]), .CK(clk), .Q(out[61])
         );
  SDFF_X1 out_reg_62_ ( .D(1'b0), .SI(n65), .SE(in[62]), .CK(clk), .Q(out[62])
         );
  INV_X2 U3 ( .A(reset), .ZN(n65) );
  AND2_X1 U67 ( .A1(in[63]), .A2(n65), .ZN(n64) );
endmodule


module regN_N32_1 ( clk, reset, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, reset;
  wire   n1, n2, n3, n5, n10, n34, n35, n36, n37;

  SDFF_X1 out_reg_31_ ( .D(1'b0), .SI(n34), .SE(in[31]), .CK(clk), .Q(out[31])
         );
  SDFF_X1 out_reg_30_ ( .D(1'b0), .SI(n34), .SE(in[30]), .CK(clk), .Q(out[30])
         );
  SDFF_X1 out_reg_29_ ( .D(1'b0), .SI(n34), .SE(in[29]), .CK(clk), .Q(out[29])
         );
  SDFF_X1 out_reg_28_ ( .D(1'b0), .SI(n34), .SE(in[28]), .CK(clk), .Q(out[28])
         );
  SDFF_X1 out_reg_27_ ( .D(1'b0), .SI(n34), .SE(in[27]), .CK(clk), .Q(out[27])
         );
  SDFF_X1 out_reg_26_ ( .D(1'b0), .SI(n34), .SE(in[26]), .CK(clk), .Q(out[26])
         );
  SDFF_X1 out_reg_25_ ( .D(1'b0), .SI(n34), .SE(in[25]), .CK(clk), .Q(out[25])
         );
  SDFF_X1 out_reg_24_ ( .D(1'b0), .SI(n34), .SE(in[24]), .CK(clk), .Q(out[24])
         );
  SDFF_X1 out_reg_23_ ( .D(1'b0), .SI(n34), .SE(in[23]), .CK(clk), .Q(out[23])
         );
  SDFF_X1 out_reg_22_ ( .D(1'b0), .SI(n34), .SE(in[22]), .CK(clk), .Q(out[22])
         );
  SDFF_X1 out_reg_21_ ( .D(1'b0), .SI(n34), .SE(in[21]), .CK(clk), .Q(out[21])
         );
  SDFF_X1 out_reg_20_ ( .D(1'b0), .SI(n35), .SE(in[20]), .CK(clk), .Q(out[20])
         );
  SDFF_X1 out_reg_19_ ( .D(1'b0), .SI(n35), .SE(in[19]), .CK(clk), .Q(out[19])
         );
  SDFF_X1 out_reg_18_ ( .D(1'b0), .SI(n35), .SE(in[18]), .CK(clk), .Q(out[18])
         );
  SDFF_X1 out_reg_17_ ( .D(1'b0), .SI(n35), .SE(in[17]), .CK(clk), .Q(out[17])
         );
  SDFF_X1 out_reg_16_ ( .D(1'b0), .SI(n35), .SE(in[16]), .CK(clk), .Q(out[16])
         );
  SDFF_X1 out_reg_15_ ( .D(1'b0), .SI(n35), .SE(in[15]), .CK(clk), .Q(out[15])
         );
  SDFF_X1 out_reg_14_ ( .D(1'b0), .SI(n35), .SE(in[14]), .CK(clk), .Q(out[14])
         );
  SDFF_X1 out_reg_13_ ( .D(1'b0), .SI(n35), .SE(in[13]), .CK(clk), .Q(out[13])
         );
  SDFF_X1 out_reg_12_ ( .D(1'b0), .SI(n35), .SE(in[12]), .CK(clk), .Q(out[12])
         );
  SDFF_X1 out_reg_11_ ( .D(1'b0), .SI(n35), .SE(in[11]), .CK(clk), .Q(out[11])
         );
  SDFF_X1 out_reg_10_ ( .D(1'b0), .SI(n35), .SE(in[10]), .CK(clk), .Q(out[10])
         );
  SDFF_X1 out_reg_8_ ( .D(1'b0), .SI(n36), .SE(in[8]), .CK(clk), .Q(out[8]) );
  SDFF_X1 out_reg_7_ ( .D(1'b0), .SI(n36), .SE(in[7]), .CK(clk), .Q(out[7]) );
  SDFF_X1 out_reg_6_ ( .D(1'b0), .SI(n36), .SE(in[6]), .CK(clk), .Q(out[6]) );
  SDFF_X1 out_reg_5_ ( .D(1'b0), .SI(n36), .SE(in[5]), .CK(clk), .Q(out[5]) );
  SDFF_X1 out_reg_3_ ( .D(1'b0), .SI(n36), .SE(in[3]), .CK(clk), .Q(out[3]) );
  DFF_X1 out_reg_2_ ( .D(n10), .CK(clk), .Q(out[2]) );
  DFF_X1 out_reg_0_ ( .D(n5), .CK(clk), .Q(out[0]) );
  DFF_X1 out_reg_1_ ( .D(n3), .CK(clk), .Q(out[1]) );
  DFF_X1 out_reg_4_ ( .D(n2), .CK(clk), .Q(out[4]) );
  DFF_X1 out_reg_9_ ( .D(n1), .CK(clk), .Q(out[9]) );
  AND2_X1 U3 ( .A1(in[9]), .A2(n36), .ZN(n1) );
  BUF_X1 U4 ( .A(n37), .Z(n35) );
  BUF_X1 U5 ( .A(n37), .Z(n34) );
  BUF_X1 U7 ( .A(n37), .Z(n36) );
  INV_X1 U12 ( .A(reset), .ZN(n37) );
  AND2_X1 U35 ( .A1(in[4]), .A2(n36), .ZN(n2) );
  AND2_X1 U36 ( .A1(in[1]), .A2(n36), .ZN(n3) );
  AND2_X1 U37 ( .A1(in[0]), .A2(n36), .ZN(n5) );
  AND2_X1 U38 ( .A1(in[2]), .A2(n36), .ZN(n10) );
endmodule


module TMSeq ( A, B, clk, reset, result );
  input [31:0] A;
  input [31:0] B;
  output [63:0] result;
  input clk, reset;

  wire   [31:0] AReg;
  wire   [31:0] BReg;
  wire   [63:0] resultReg;

  regN_N32_0 regA ( .clk(clk), .reset(reset), .in(A), .out(AReg) );
  regN_N32_1 regB ( .clk(clk), .reset(reset), .in(B), .out(BReg) );
  TM multiplier ( .a(AReg), .b(BReg), .result(resultReg) );
  regN_N64 outA ( .clk(clk), .reset(reset), .in(resultReg), .out(result) );
endmodule



module FullAdder_0 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_3 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_4 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_5 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_6 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_7 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_8 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_9 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_10 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_11 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_12 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_13 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_14 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_15 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_16 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_17 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_18 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_19 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_20 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_21 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_22 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_23 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_24 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_25 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_26 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_27 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_28 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_29 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_30 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_31 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder ( a, b, cin, sum, cout, overflow );
  input [31:0] a;
  input [31:0] b;
  output [31:0] sum;
  input cin;
  output cout, overflow;
  wire   n3, n4;
  wire   [30:0] passCout;

  FullAdder_0 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_31 bit1 ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(sum[1]), 
        .cout(passCout[1]) );
  FullAdder_30 bit2 ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(sum[2]), 
        .cout(passCout[2]) );
  FullAdder_29 bit3 ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(sum[3]), 
        .cout(passCout[3]) );
  FullAdder_28 bit4 ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(sum[4]), 
        .cout(passCout[4]) );
  FullAdder_27 bit5 ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(sum[5]), 
        .cout(passCout[5]) );
  FullAdder_26 bit6 ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(sum[6]), 
        .cout(passCout[6]) );
  FullAdder_25 bit7 ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(sum[7]), 
        .cout(passCout[7]) );
  FullAdder_24 bit8 ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(sum[8]), 
        .cout(passCout[8]) );
  FullAdder_23 bit9 ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(sum[9]), 
        .cout(passCout[9]) );
  FullAdder_22 bit10 ( .a(a[10]), .b(b[10]), .cin(passCout[9]), .sum(sum[10]), 
        .cout(passCout[10]) );
  FullAdder_21 bit11 ( .a(a[11]), .b(b[11]), .cin(passCout[10]), .sum(sum[11]), 
        .cout(passCout[11]) );
  FullAdder_20 bit12 ( .a(a[12]), .b(b[12]), .cin(passCout[11]), .sum(sum[12]), 
        .cout(passCout[12]) );
  FullAdder_19 bit13 ( .a(a[13]), .b(b[13]), .cin(passCout[12]), .sum(sum[13]), 
        .cout(passCout[13]) );
  FullAdder_18 bit14 ( .a(a[14]), .b(b[14]), .cin(passCout[13]), .sum(sum[14]), 
        .cout(passCout[14]) );
  FullAdder_17 bit15 ( .a(a[15]), .b(b[15]), .cin(passCout[14]), .sum(sum[15]), 
        .cout(passCout[15]) );
  FullAdder_16 bit16 ( .a(a[16]), .b(b[16]), .cin(passCout[15]), .sum(sum[16]), 
        .cout(passCout[16]) );
  FullAdder_15 bit17 ( .a(a[17]), .b(b[17]), .cin(passCout[16]), .sum(sum[17]), 
        .cout(passCout[17]) );
  FullAdder_14 bit18 ( .a(a[18]), .b(b[18]), .cin(passCout[17]), .sum(sum[18]), 
        .cout(passCout[18]) );
  FullAdder_13 bit19 ( .a(a[19]), .b(b[19]), .cin(passCout[18]), .sum(sum[19]), 
        .cout(passCout[19]) );
  FullAdder_12 bit20 ( .a(a[20]), .b(b[20]), .cin(passCout[19]), .sum(sum[20]), 
        .cout(passCout[20]) );
  FullAdder_11 bit21 ( .a(a[21]), .b(b[21]), .cin(passCout[20]), .sum(sum[21]), 
        .cout(passCout[21]) );
  FullAdder_10 bit22 ( .a(a[22]), .b(b[22]), .cin(passCout[21]), .sum(sum[22]), 
        .cout(passCout[22]) );
  FullAdder_9 bit23 ( .a(a[23]), .b(b[23]), .cin(passCout[22]), .sum(sum[23]), 
        .cout(passCout[23]) );
  FullAdder_8 bit24 ( .a(a[24]), .b(b[24]), .cin(passCout[23]), .sum(sum[24]), 
        .cout(passCout[24]) );
  FullAdder_7 bit25 ( .a(a[25]), .b(b[25]), .cin(passCout[24]), .sum(sum[25]), 
        .cout(passCout[25]) );
  FullAdder_6 bit26 ( .a(a[26]), .b(b[26]), .cin(passCout[25]), .sum(sum[26]), 
        .cout(passCout[26]) );
  FullAdder_5 bit27 ( .a(a[27]), .b(b[27]), .cin(passCout[26]), .sum(sum[27]), 
        .cout(passCout[27]) );
  FullAdder_4 bit28 ( .a(a[28]), .b(b[28]), .cin(passCout[27]), .sum(sum[28]), 
        .cout(passCout[28]) );
  FullAdder_3 bit29 ( .a(a[29]), .b(b[29]), .cin(passCout[28]), .sum(sum[29]), 
        .cout(passCout[29]) );
  FullAdder_2 bit30 ( .a(a[30]), .b(b[30]), .cin(passCout[29]), .sum(sum[30]), 
        .cout(passCout[30]) );
  FullAdder_1 bit31 ( .a(a[31]), .b(b[31]), .cin(passCout[30]), .sum(sum[31]), 
        .cout(cout) );
  NOR2_X1 U4 ( .A1(n3), .A2(n4), .ZN(overflow) );
  XOR2_X1 U5 ( .A(b[31]), .B(a[31]), .Z(n4) );
  XNOR2_X1 U6 ( .A(a[31]), .B(sum[31]), .ZN(n3) );
endmodule


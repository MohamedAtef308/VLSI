
module regN_N32_0 ( clk, reset, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, reset;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  DFF_X1 out_reg_9_ ( .D(n32), .CK(clk), .Q(out[9]) );
  DFF_X1 out_reg_8_ ( .D(n31), .CK(clk), .Q(out[8]) );
  DFF_X1 out_reg_7_ ( .D(n30), .CK(clk), .Q(out[7]) );
  DFF_X1 out_reg_6_ ( .D(n29), .CK(clk), .Q(out[6]) );
  DFF_X1 out_reg_5_ ( .D(n28), .CK(clk), .Q(out[5]) );
  DFF_X1 out_reg_4_ ( .D(n27), .CK(clk), .Q(out[4]) );
  DFF_X1 out_reg_3_ ( .D(n26), .CK(clk), .Q(out[3]) );
  DFF_X1 out_reg_2_ ( .D(n25), .CK(clk), .Q(out[2]) );
  DFF_X1 out_reg_1_ ( .D(n24), .CK(clk), .Q(out[1]) );
  DFF_X1 out_reg_0_ ( .D(n23), .CK(clk), .Q(out[0]) );
  DFF_X1 out_reg_31_ ( .D(n22), .CK(clk), .Q(out[31]) );
  DFF_X1 out_reg_30_ ( .D(n21), .CK(clk), .Q(out[30]) );
  DFF_X1 out_reg_29_ ( .D(n20), .CK(clk), .Q(out[29]) );
  DFF_X1 out_reg_28_ ( .D(n19), .CK(clk), .Q(out[28]) );
  DFF_X1 out_reg_27_ ( .D(n18), .CK(clk), .Q(out[27]) );
  DFF_X1 out_reg_26_ ( .D(n17), .CK(clk), .Q(out[26]) );
  DFF_X1 out_reg_25_ ( .D(n16), .CK(clk), .Q(out[25]) );
  DFF_X1 out_reg_24_ ( .D(n15), .CK(clk), .Q(out[24]) );
  DFF_X1 out_reg_23_ ( .D(n14), .CK(clk), .Q(out[23]) );
  DFF_X1 out_reg_22_ ( .D(n13), .CK(clk), .Q(out[22]) );
  DFF_X1 out_reg_21_ ( .D(n12), .CK(clk), .Q(out[21]) );
  DFF_X1 out_reg_20_ ( .D(n11), .CK(clk), .Q(out[20]) );
  DFF_X1 out_reg_19_ ( .D(n10), .CK(clk), .Q(out[19]) );
  DFF_X1 out_reg_18_ ( .D(n9), .CK(clk), .Q(out[18]) );
  DFF_X1 out_reg_17_ ( .D(n8), .CK(clk), .Q(out[17]) );
  DFF_X1 out_reg_16_ ( .D(n7), .CK(clk), .Q(out[16]) );
  DFF_X1 out_reg_15_ ( .D(n6), .CK(clk), .Q(out[15]) );
  DFF_X1 out_reg_14_ ( .D(n5), .CK(clk), .Q(out[14]) );
  DFF_X1 out_reg_13_ ( .D(n4), .CK(clk), .Q(out[13]) );
  DFF_X1 out_reg_12_ ( .D(n3), .CK(clk), .Q(out[12]) );
  DFF_X1 out_reg_11_ ( .D(n2), .CK(clk), .Q(out[11]) );
  DFF_X1 out_reg_10_ ( .D(n1), .CK(clk), .Q(out[10]) );
  AND2_X1 U3 ( .A1(in[10]), .A2(n34), .ZN(n1) );
  AND2_X1 U4 ( .A1(in[11]), .A2(n34), .ZN(n2) );
  AND2_X1 U5 ( .A1(in[12]), .A2(n34), .ZN(n3) );
  AND2_X1 U6 ( .A1(in[13]), .A2(n34), .ZN(n4) );
  AND2_X1 U7 ( .A1(in[14]), .A2(n34), .ZN(n5) );
  AND2_X1 U8 ( .A1(in[15]), .A2(n34), .ZN(n6) );
  AND2_X1 U9 ( .A1(in[16]), .A2(n34), .ZN(n7) );
  AND2_X1 U10 ( .A1(in[17]), .A2(n34), .ZN(n8) );
  AND2_X1 U11 ( .A1(in[18]), .A2(n34), .ZN(n9) );
  AND2_X1 U12 ( .A1(in[19]), .A2(n34), .ZN(n10) );
  AND2_X1 U13 ( .A1(in[20]), .A2(n34), .ZN(n11) );
  AND2_X1 U14 ( .A1(in[21]), .A2(n33), .ZN(n12) );
  AND2_X1 U15 ( .A1(in[22]), .A2(n33), .ZN(n13) );
  AND2_X1 U16 ( .A1(in[23]), .A2(n33), .ZN(n14) );
  AND2_X1 U17 ( .A1(in[24]), .A2(n33), .ZN(n15) );
  AND2_X1 U18 ( .A1(in[25]), .A2(n33), .ZN(n16) );
  AND2_X1 U19 ( .A1(in[26]), .A2(n33), .ZN(n17) );
  AND2_X1 U20 ( .A1(in[27]), .A2(n33), .ZN(n18) );
  AND2_X1 U21 ( .A1(in[28]), .A2(n33), .ZN(n19) );
  AND2_X1 U22 ( .A1(in[29]), .A2(n33), .ZN(n20) );
  AND2_X1 U23 ( .A1(in[30]), .A2(n33), .ZN(n21) );
  AND2_X1 U24 ( .A1(in[31]), .A2(n33), .ZN(n22) );
  AND2_X1 U25 ( .A1(in[0]), .A2(n35), .ZN(n23) );
  AND2_X1 U26 ( .A1(in[1]), .A2(n35), .ZN(n24) );
  AND2_X1 U27 ( .A1(in[2]), .A2(n35), .ZN(n25) );
  AND2_X1 U28 ( .A1(in[3]), .A2(n35), .ZN(n26) );
  AND2_X1 U29 ( .A1(in[4]), .A2(n35), .ZN(n27) );
  AND2_X1 U30 ( .A1(in[5]), .A2(n35), .ZN(n28) );
  AND2_X1 U31 ( .A1(in[6]), .A2(n35), .ZN(n29) );
  AND2_X1 U32 ( .A1(in[7]), .A2(n35), .ZN(n30) );
  AND2_X1 U33 ( .A1(in[8]), .A2(n35), .ZN(n31) );
  AND2_X1 U34 ( .A1(in[9]), .A2(n35), .ZN(n32) );
  BUF_X1 U35 ( .A(n36), .Z(n34) );
  BUF_X1 U36 ( .A(n36), .Z(n33) );
  INV_X1 U37 ( .A(reset), .ZN(n36) );
  BUF_X1 U38 ( .A(n36), .Z(n35) );
endmodule


module regN_N32_2 ( clk, reset, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, reset;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  DFF_X1 out_reg_9_ ( .D(n32), .CK(clk), .Q(out[9]) );
  DFF_X1 out_reg_8_ ( .D(n31), .CK(clk), .Q(out[8]) );
  DFF_X1 out_reg_7_ ( .D(n30), .CK(clk), .Q(out[7]) );
  DFF_X1 out_reg_6_ ( .D(n29), .CK(clk), .Q(out[6]) );
  DFF_X1 out_reg_5_ ( .D(n28), .CK(clk), .Q(out[5]) );
  DFF_X1 out_reg_4_ ( .D(n27), .CK(clk), .Q(out[4]) );
  DFF_X1 out_reg_3_ ( .D(n26), .CK(clk), .Q(out[3]) );
  DFF_X1 out_reg_2_ ( .D(n25), .CK(clk), .Q(out[2]) );
  DFF_X1 out_reg_1_ ( .D(n24), .CK(clk), .Q(out[1]) );
  DFF_X1 out_reg_0_ ( .D(n23), .CK(clk), .Q(out[0]) );
  DFF_X1 out_reg_31_ ( .D(n22), .CK(clk), .Q(out[31]) );
  DFF_X1 out_reg_30_ ( .D(n21), .CK(clk), .Q(out[30]) );
  DFF_X1 out_reg_29_ ( .D(n20), .CK(clk), .Q(out[29]) );
  DFF_X1 out_reg_28_ ( .D(n19), .CK(clk), .Q(out[28]) );
  DFF_X1 out_reg_27_ ( .D(n18), .CK(clk), .Q(out[27]) );
  DFF_X1 out_reg_26_ ( .D(n17), .CK(clk), .Q(out[26]) );
  DFF_X1 out_reg_25_ ( .D(n16), .CK(clk), .Q(out[25]) );
  DFF_X1 out_reg_24_ ( .D(n15), .CK(clk), .Q(out[24]) );
  DFF_X1 out_reg_23_ ( .D(n14), .CK(clk), .Q(out[23]) );
  DFF_X1 out_reg_22_ ( .D(n13), .CK(clk), .Q(out[22]) );
  DFF_X1 out_reg_21_ ( .D(n12), .CK(clk), .Q(out[21]) );
  DFF_X1 out_reg_20_ ( .D(n11), .CK(clk), .Q(out[20]) );
  DFF_X1 out_reg_19_ ( .D(n10), .CK(clk), .Q(out[19]) );
  DFF_X1 out_reg_18_ ( .D(n9), .CK(clk), .Q(out[18]) );
  DFF_X1 out_reg_17_ ( .D(n8), .CK(clk), .Q(out[17]) );
  DFF_X1 out_reg_16_ ( .D(n7), .CK(clk), .Q(out[16]) );
  DFF_X1 out_reg_15_ ( .D(n6), .CK(clk), .Q(out[15]) );
  DFF_X1 out_reg_14_ ( .D(n5), .CK(clk), .Q(out[14]) );
  DFF_X1 out_reg_13_ ( .D(n4), .CK(clk), .Q(out[13]) );
  DFF_X1 out_reg_12_ ( .D(n3), .CK(clk), .Q(out[12]) );
  DFF_X1 out_reg_11_ ( .D(n2), .CK(clk), .Q(out[11]) );
  DFF_X1 out_reg_10_ ( .D(n1), .CK(clk), .Q(out[10]) );
  AND2_X1 U3 ( .A1(in[10]), .A2(n34), .ZN(n1) );
  AND2_X1 U4 ( .A1(in[11]), .A2(n34), .ZN(n2) );
  AND2_X1 U5 ( .A1(in[12]), .A2(n34), .ZN(n3) );
  AND2_X1 U6 ( .A1(in[13]), .A2(n34), .ZN(n4) );
  AND2_X1 U7 ( .A1(in[14]), .A2(n34), .ZN(n5) );
  AND2_X1 U8 ( .A1(in[15]), .A2(n34), .ZN(n6) );
  AND2_X1 U9 ( .A1(in[16]), .A2(n34), .ZN(n7) );
  AND2_X1 U10 ( .A1(in[17]), .A2(n34), .ZN(n8) );
  AND2_X1 U11 ( .A1(in[18]), .A2(n34), .ZN(n9) );
  AND2_X1 U12 ( .A1(in[19]), .A2(n34), .ZN(n10) );
  AND2_X1 U13 ( .A1(in[20]), .A2(n34), .ZN(n11) );
  AND2_X1 U14 ( .A1(in[21]), .A2(n33), .ZN(n12) );
  AND2_X1 U15 ( .A1(in[22]), .A2(n33), .ZN(n13) );
  AND2_X1 U16 ( .A1(in[23]), .A2(n33), .ZN(n14) );
  AND2_X1 U17 ( .A1(in[24]), .A2(n33), .ZN(n15) );
  AND2_X1 U18 ( .A1(in[25]), .A2(n33), .ZN(n16) );
  AND2_X1 U19 ( .A1(in[26]), .A2(n33), .ZN(n17) );
  AND2_X1 U20 ( .A1(in[27]), .A2(n33), .ZN(n18) );
  AND2_X1 U21 ( .A1(in[28]), .A2(n33), .ZN(n19) );
  AND2_X1 U22 ( .A1(in[29]), .A2(n33), .ZN(n20) );
  AND2_X1 U23 ( .A1(in[30]), .A2(n33), .ZN(n21) );
  AND2_X1 U24 ( .A1(in[31]), .A2(n33), .ZN(n22) );
  AND2_X1 U25 ( .A1(in[0]), .A2(n35), .ZN(n23) );
  AND2_X1 U26 ( .A1(in[1]), .A2(n35), .ZN(n24) );
  AND2_X1 U27 ( .A1(in[2]), .A2(n35), .ZN(n25) );
  AND2_X1 U28 ( .A1(in[3]), .A2(n35), .ZN(n26) );
  AND2_X1 U29 ( .A1(in[4]), .A2(n35), .ZN(n27) );
  AND2_X1 U30 ( .A1(in[5]), .A2(n35), .ZN(n28) );
  AND2_X1 U31 ( .A1(in[6]), .A2(n35), .ZN(n29) );
  AND2_X1 U32 ( .A1(in[7]), .A2(n35), .ZN(n30) );
  AND2_X1 U33 ( .A1(in[8]), .A2(n35), .ZN(n31) );
  AND2_X1 U34 ( .A1(in[9]), .A2(n35), .ZN(n32) );
  BUF_X1 U35 ( .A(n36), .Z(n35) );
  INV_X1 U36 ( .A(reset), .ZN(n36) );
  BUF_X1 U37 ( .A(n36), .Z(n34) );
  BUF_X1 U38 ( .A(n36), .Z(n33) );
endmodule


module FPM_DW01_add_2 ( A, B, CI, SUM, CO );
  input [45:0] A;
  input [45:0] B;
  output [45:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110;
  assign SUM[22] = A[22];
  assign SUM[21] = A[21];

  AND2_X1 U2 ( .A1(n2), .A2(n110), .ZN(SUM[23]) );
  INV_X1 U3 ( .A(n93), .ZN(n21) );
  INV_X1 U4 ( .A(n85), .ZN(n19) );
  INV_X1 U5 ( .A(n69), .ZN(n15) );
  INV_X1 U6 ( .A(n61), .ZN(n13) );
  INV_X1 U7 ( .A(n53), .ZN(n11) );
  INV_X1 U8 ( .A(n45), .ZN(n9) );
  INV_X1 U9 ( .A(n37), .ZN(n7) );
  INV_X1 U10 ( .A(n77), .ZN(n17) );
  INV_X1 U11 ( .A(n55), .ZN(n12) );
  INV_X1 U12 ( .A(n47), .ZN(n10) );
  INV_X1 U13 ( .A(n39), .ZN(n8) );
  INV_X1 U14 ( .A(n31), .ZN(n6) );
  INV_X1 U15 ( .A(n101), .ZN(n23) );
  INV_X1 U16 ( .A(n103), .ZN(n24) );
  INV_X1 U17 ( .A(n87), .ZN(n20) );
  INV_X1 U18 ( .A(n79), .ZN(n18) );
  INV_X1 U19 ( .A(n63), .ZN(n14) );
  INV_X1 U20 ( .A(n95), .ZN(n22) );
  INV_X1 U21 ( .A(n71), .ZN(n16) );
  INV_X1 U22 ( .A(n4), .ZN(n110) );
  INV_X1 U23 ( .A(n29), .ZN(n5) );
  AND2_X1 U24 ( .A1(B[23]), .A2(A[23]), .ZN(n4) );
  OR2_X1 U25 ( .A1(B[23]), .A2(A[23]), .ZN(n2) );
  AOI21_X1 U26 ( .B1(n99), .B2(n23), .A(n100), .ZN(n3) );
  XOR2_X1 U27 ( .A(A[44]), .B(n26), .Z(SUM[45]) );
  INV_X1 U28 ( .A(n108), .ZN(n25) );
  AOI21_X1 U29 ( .B1(n27), .B2(n5), .A(n28), .ZN(n26) );
  XOR2_X1 U30 ( .A(n27), .B(n30), .Z(SUM[44]) );
  NOR2_X1 U31 ( .A1(n28), .A2(n29), .ZN(n30) );
  NOR2_X1 U32 ( .A1(B[44]), .A2(A[44]), .ZN(n29) );
  AND2_X1 U33 ( .A1(B[44]), .A2(A[44]), .ZN(n28) );
  OAI21_X1 U34 ( .B1(n31), .B2(n32), .A(n33), .ZN(n27) );
  XOR2_X1 U35 ( .A(n34), .B(n32), .Z(SUM[43]) );
  AOI21_X1 U36 ( .B1(n7), .B2(n35), .A(n36), .ZN(n32) );
  NAND2_X1 U37 ( .A1(n6), .A2(n33), .ZN(n34) );
  NAND2_X1 U38 ( .A1(B[43]), .A2(A[43]), .ZN(n33) );
  NOR2_X1 U39 ( .A1(B[43]), .A2(A[43]), .ZN(n31) );
  XOR2_X1 U40 ( .A(n35), .B(n38), .Z(SUM[42]) );
  NOR2_X1 U41 ( .A1(n36), .A2(n37), .ZN(n38) );
  NOR2_X1 U42 ( .A1(B[42]), .A2(A[42]), .ZN(n37) );
  AND2_X1 U43 ( .A1(B[42]), .A2(A[42]), .ZN(n36) );
  OAI21_X1 U44 ( .B1(n39), .B2(n40), .A(n41), .ZN(n35) );
  XOR2_X1 U45 ( .A(n42), .B(n40), .Z(SUM[41]) );
  AOI21_X1 U46 ( .B1(n9), .B2(n43), .A(n44), .ZN(n40) );
  NAND2_X1 U47 ( .A1(n8), .A2(n41), .ZN(n42) );
  NAND2_X1 U48 ( .A1(B[41]), .A2(A[41]), .ZN(n41) );
  NOR2_X1 U49 ( .A1(B[41]), .A2(A[41]), .ZN(n39) );
  XOR2_X1 U50 ( .A(n43), .B(n46), .Z(SUM[40]) );
  NOR2_X1 U51 ( .A1(n44), .A2(n45), .ZN(n46) );
  NOR2_X1 U52 ( .A1(B[40]), .A2(A[40]), .ZN(n45) );
  AND2_X1 U53 ( .A1(B[40]), .A2(A[40]), .ZN(n44) );
  OAI21_X1 U54 ( .B1(n47), .B2(n48), .A(n49), .ZN(n43) );
  XOR2_X1 U55 ( .A(n50), .B(n48), .Z(SUM[39]) );
  AOI21_X1 U56 ( .B1(n11), .B2(n51), .A(n52), .ZN(n48) );
  NAND2_X1 U57 ( .A1(n10), .A2(n49), .ZN(n50) );
  NAND2_X1 U58 ( .A1(B[39]), .A2(A[39]), .ZN(n49) );
  NOR2_X1 U59 ( .A1(B[39]), .A2(A[39]), .ZN(n47) );
  XOR2_X1 U60 ( .A(n51), .B(n54), .Z(SUM[38]) );
  NOR2_X1 U61 ( .A1(n52), .A2(n53), .ZN(n54) );
  NOR2_X1 U62 ( .A1(B[38]), .A2(A[38]), .ZN(n53) );
  AND2_X1 U63 ( .A1(B[38]), .A2(A[38]), .ZN(n52) );
  OAI21_X1 U64 ( .B1(n55), .B2(n56), .A(n57), .ZN(n51) );
  XOR2_X1 U65 ( .A(n58), .B(n56), .Z(SUM[37]) );
  AOI21_X1 U66 ( .B1(n13), .B2(n59), .A(n60), .ZN(n56) );
  NAND2_X1 U67 ( .A1(n12), .A2(n57), .ZN(n58) );
  NAND2_X1 U68 ( .A1(B[37]), .A2(A[37]), .ZN(n57) );
  NOR2_X1 U69 ( .A1(B[37]), .A2(A[37]), .ZN(n55) );
  XOR2_X1 U70 ( .A(n59), .B(n62), .Z(SUM[36]) );
  NOR2_X1 U71 ( .A1(n60), .A2(n61), .ZN(n62) );
  NOR2_X1 U72 ( .A1(B[36]), .A2(A[36]), .ZN(n61) );
  AND2_X1 U73 ( .A1(B[36]), .A2(A[36]), .ZN(n60) );
  OAI21_X1 U74 ( .B1(n63), .B2(n64), .A(n65), .ZN(n59) );
  XOR2_X1 U75 ( .A(n66), .B(n64), .Z(SUM[35]) );
  AOI21_X1 U76 ( .B1(n15), .B2(n67), .A(n68), .ZN(n64) );
  NAND2_X1 U77 ( .A1(n14), .A2(n65), .ZN(n66) );
  NAND2_X1 U78 ( .A1(B[35]), .A2(A[35]), .ZN(n65) );
  NOR2_X1 U79 ( .A1(B[35]), .A2(A[35]), .ZN(n63) );
  XOR2_X1 U80 ( .A(n67), .B(n70), .Z(SUM[34]) );
  NOR2_X1 U81 ( .A1(n68), .A2(n69), .ZN(n70) );
  NOR2_X1 U82 ( .A1(B[34]), .A2(A[34]), .ZN(n69) );
  AND2_X1 U83 ( .A1(B[34]), .A2(A[34]), .ZN(n68) );
  OAI21_X1 U84 ( .B1(n71), .B2(n72), .A(n73), .ZN(n67) );
  XOR2_X1 U85 ( .A(n74), .B(n72), .Z(SUM[33]) );
  AOI21_X1 U86 ( .B1(n17), .B2(n75), .A(n76), .ZN(n72) );
  NAND2_X1 U87 ( .A1(n16), .A2(n73), .ZN(n74) );
  NAND2_X1 U88 ( .A1(B[33]), .A2(A[33]), .ZN(n73) );
  NOR2_X1 U89 ( .A1(B[33]), .A2(A[33]), .ZN(n71) );
  XOR2_X1 U90 ( .A(n75), .B(n78), .Z(SUM[32]) );
  NOR2_X1 U91 ( .A1(n76), .A2(n77), .ZN(n78) );
  NOR2_X1 U92 ( .A1(B[32]), .A2(A[32]), .ZN(n77) );
  AND2_X1 U93 ( .A1(B[32]), .A2(A[32]), .ZN(n76) );
  OAI21_X1 U94 ( .B1(n79), .B2(n80), .A(n81), .ZN(n75) );
  XOR2_X1 U95 ( .A(n82), .B(n80), .Z(SUM[31]) );
  AOI21_X1 U96 ( .B1(n19), .B2(n83), .A(n84), .ZN(n80) );
  NAND2_X1 U97 ( .A1(n18), .A2(n81), .ZN(n82) );
  NAND2_X1 U98 ( .A1(B[31]), .A2(A[31]), .ZN(n81) );
  NOR2_X1 U99 ( .A1(B[31]), .A2(A[31]), .ZN(n79) );
  XOR2_X1 U100 ( .A(n83), .B(n86), .Z(SUM[30]) );
  NOR2_X1 U101 ( .A1(n84), .A2(n85), .ZN(n86) );
  NOR2_X1 U102 ( .A1(B[30]), .A2(A[30]), .ZN(n85) );
  AND2_X1 U103 ( .A1(B[30]), .A2(A[30]), .ZN(n84) );
  OAI21_X1 U104 ( .B1(n87), .B2(n88), .A(n89), .ZN(n83) );
  XOR2_X1 U105 ( .A(n90), .B(n88), .Z(SUM[29]) );
  AOI21_X1 U106 ( .B1(n21), .B2(n91), .A(n92), .ZN(n88) );
  NAND2_X1 U107 ( .A1(n20), .A2(n89), .ZN(n90) );
  NAND2_X1 U108 ( .A1(B[29]), .A2(A[29]), .ZN(n89) );
  NOR2_X1 U109 ( .A1(B[29]), .A2(A[29]), .ZN(n87) );
  XOR2_X1 U110 ( .A(n91), .B(n94), .Z(SUM[28]) );
  NOR2_X1 U111 ( .A1(n92), .A2(n93), .ZN(n94) );
  NOR2_X1 U112 ( .A1(B[28]), .A2(A[28]), .ZN(n93) );
  AND2_X1 U113 ( .A1(B[28]), .A2(A[28]), .ZN(n92) );
  OAI21_X1 U114 ( .B1(n95), .B2(n96), .A(n97), .ZN(n91) );
  XOR2_X1 U115 ( .A(n98), .B(n3), .Z(SUM[27]) );
  AOI21_X1 U116 ( .B1(n99), .B2(n23), .A(n100), .ZN(n96) );
  NAND2_X1 U117 ( .A1(n22), .A2(n97), .ZN(n98) );
  NAND2_X1 U118 ( .A1(B[27]), .A2(A[27]), .ZN(n97) );
  NOR2_X1 U119 ( .A1(B[27]), .A2(A[27]), .ZN(n95) );
  XOR2_X1 U120 ( .A(n99), .B(n102), .Z(SUM[26]) );
  NOR2_X1 U121 ( .A1(n100), .A2(n101), .ZN(n102) );
  NOR2_X1 U122 ( .A1(B[26]), .A2(A[26]), .ZN(n101) );
  AND2_X1 U123 ( .A1(B[26]), .A2(A[26]), .ZN(n100) );
  OAI21_X1 U124 ( .B1(n103), .B2(n104), .A(n105), .ZN(n99) );
  XOR2_X1 U125 ( .A(n106), .B(n104), .Z(SUM[25]) );
  AOI21_X1 U126 ( .B1(n25), .B2(n4), .A(n107), .ZN(n104) );
  NAND2_X1 U127 ( .A1(n24), .A2(n105), .ZN(n106) );
  NAND2_X1 U128 ( .A1(B[25]), .A2(A[25]), .ZN(n105) );
  NOR2_X1 U129 ( .A1(B[25]), .A2(A[25]), .ZN(n103) );
  XOR2_X1 U130 ( .A(n4), .B(n109), .Z(SUM[24]) );
  NOR2_X1 U131 ( .A1(n107), .A2(n108), .ZN(n109) );
  NOR2_X1 U132 ( .A1(B[24]), .A2(A[24]), .ZN(n108) );
  AND2_X1 U133 ( .A1(B[24]), .A2(A[24]), .ZN(n107) );
endmodule


module FPM_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   ab_22__22_, ab_22__21_, ab_22__20_, ab_22__19_, ab_22__18_,
         ab_22__17_, ab_22__16_, ab_22__15_, ab_22__14_, ab_22__13_,
         ab_22__12_, ab_22__11_, ab_22__10_, ab_22__9_, ab_22__8_, ab_22__7_,
         ab_22__6_, ab_22__5_, ab_22__4_, ab_22__3_, ab_22__2_, ab_22__1_,
         ab_22__0_, ab_21__22_, ab_21__21_, ab_21__20_, ab_21__19_, ab_21__18_,
         ab_21__17_, ab_21__16_, ab_21__15_, ab_21__14_, ab_21__13_,
         ab_21__12_, ab_21__11_, ab_21__10_, ab_21__9_, ab_21__8_, ab_21__7_,
         ab_21__6_, ab_21__5_, ab_21__4_, ab_21__3_, ab_21__2_, ab_21__1_,
         ab_21__0_, ab_20__22_, ab_20__21_, ab_20__20_, ab_20__19_, ab_20__18_,
         ab_20__17_, ab_20__16_, ab_20__15_, ab_20__14_, ab_20__13_,
         ab_20__12_, ab_20__11_, ab_20__10_, ab_20__9_, ab_20__8_, ab_20__7_,
         ab_20__6_, ab_20__5_, ab_20__4_, ab_20__3_, ab_20__2_, ab_20__1_,
         ab_20__0_, ab_19__22_, ab_19__21_, ab_19__20_, ab_19__19_, ab_19__18_,
         ab_19__17_, ab_19__16_, ab_19__15_, ab_19__14_, ab_19__13_,
         ab_19__12_, ab_19__11_, ab_19__10_, ab_19__9_, ab_19__8_, ab_19__7_,
         ab_19__6_, ab_19__5_, ab_19__4_, ab_19__3_, ab_19__2_, ab_19__1_,
         ab_19__0_, ab_18__22_, ab_18__21_, ab_18__20_, ab_18__19_, ab_18__18_,
         ab_18__17_, ab_18__16_, ab_18__15_, ab_18__14_, ab_18__13_,
         ab_18__12_, ab_18__11_, ab_18__10_, ab_18__9_, ab_18__8_, ab_18__7_,
         ab_18__6_, ab_18__5_, ab_18__4_, ab_18__3_, ab_18__2_, ab_18__1_,
         ab_18__0_, ab_17__22_, ab_17__21_, ab_17__20_, ab_17__19_, ab_17__18_,
         ab_17__17_, ab_17__16_, ab_17__15_, ab_17__14_, ab_17__13_,
         ab_17__12_, ab_17__11_, ab_17__10_, ab_17__9_, ab_17__8_, ab_17__7_,
         ab_17__6_, ab_17__5_, ab_17__4_, ab_17__3_, ab_17__2_, ab_17__1_,
         ab_17__0_, ab_16__22_, ab_16__21_, ab_16__20_, ab_16__19_, ab_16__18_,
         ab_16__17_, ab_16__16_, ab_16__15_, ab_16__14_, ab_16__13_,
         ab_16__12_, ab_16__11_, ab_16__10_, ab_16__9_, ab_16__8_, ab_16__7_,
         ab_16__6_, ab_16__5_, ab_16__4_, ab_16__3_, ab_16__2_, ab_16__1_,
         ab_16__0_, ab_15__22_, ab_15__21_, ab_15__20_, ab_15__19_, ab_15__18_,
         ab_15__17_, ab_15__16_, ab_15__15_, ab_15__14_, ab_15__13_,
         ab_15__12_, ab_15__11_, ab_15__10_, ab_15__9_, ab_15__8_, ab_15__7_,
         ab_15__6_, ab_15__5_, ab_15__4_, ab_15__3_, ab_15__2_, ab_15__1_,
         ab_15__0_, ab_14__22_, ab_14__21_, ab_14__20_, ab_14__19_, ab_14__18_,
         ab_14__17_, ab_14__16_, ab_14__15_, ab_14__14_, ab_14__13_,
         ab_14__12_, ab_14__11_, ab_14__10_, ab_14__9_, ab_14__8_, ab_14__7_,
         ab_14__6_, ab_14__5_, ab_14__4_, ab_14__3_, ab_14__2_, ab_14__1_,
         ab_14__0_, ab_13__22_, ab_13__21_, ab_13__20_, ab_13__19_, ab_13__18_,
         ab_13__17_, ab_13__16_, ab_13__15_, ab_13__14_, ab_13__13_,
         ab_13__12_, ab_13__11_, ab_13__10_, ab_13__9_, ab_13__8_, ab_13__7_,
         ab_13__6_, ab_13__5_, ab_13__4_, ab_13__3_, ab_13__2_, ab_13__1_,
         ab_13__0_, ab_12__22_, ab_12__21_, ab_12__20_, ab_12__19_, ab_12__18_,
         ab_12__17_, ab_12__16_, ab_12__15_, ab_12__14_, ab_12__13_,
         ab_12__12_, ab_12__11_, ab_12__10_, ab_12__9_, ab_12__8_, ab_12__7_,
         ab_12__6_, ab_12__5_, ab_12__4_, ab_12__3_, ab_12__2_, ab_12__1_,
         ab_12__0_, ab_11__22_, ab_11__21_, ab_11__20_, ab_11__19_, ab_11__18_,
         ab_11__17_, ab_11__16_, ab_11__15_, ab_11__14_, ab_11__13_,
         ab_11__12_, ab_11__11_, ab_11__10_, ab_11__9_, ab_11__8_, ab_11__7_,
         ab_11__6_, ab_11__5_, ab_11__4_, ab_11__3_, ab_11__2_, ab_11__1_,
         ab_11__0_, ab_10__22_, ab_10__21_, ab_10__20_, ab_10__19_, ab_10__18_,
         ab_10__17_, ab_10__16_, ab_10__15_, ab_10__14_, ab_10__13_,
         ab_10__12_, ab_10__11_, ab_10__10_, ab_10__9_, ab_10__8_, ab_10__7_,
         ab_10__6_, ab_10__5_, ab_10__4_, ab_10__3_, ab_10__2_, ab_10__1_,
         ab_10__0_, ab_9__22_, ab_9__21_, ab_9__20_, ab_9__19_, ab_9__18_,
         ab_9__17_, ab_9__16_, ab_9__15_, ab_9__14_, ab_9__13_, ab_9__12_,
         ab_9__11_, ab_9__10_, ab_9__9_, ab_9__8_, ab_9__7_, ab_9__6_,
         ab_9__5_, ab_9__4_, ab_9__3_, ab_9__2_, ab_9__1_, ab_9__0_, ab_8__22_,
         ab_8__21_, ab_8__20_, ab_8__19_, ab_8__18_, ab_8__17_, ab_8__16_,
         ab_8__15_, ab_8__14_, ab_8__13_, ab_8__12_, ab_8__11_, ab_8__10_,
         ab_8__9_, ab_8__8_, ab_8__7_, ab_8__6_, ab_8__5_, ab_8__4_, ab_8__3_,
         ab_8__2_, ab_8__1_, ab_8__0_, ab_7__22_, ab_7__21_, ab_7__20_,
         ab_7__19_, ab_7__18_, ab_7__17_, ab_7__16_, ab_7__15_, ab_7__14_,
         ab_7__13_, ab_7__12_, ab_7__11_, ab_7__10_, ab_7__9_, ab_7__8_,
         ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__22_, ab_6__21_, ab_6__20_, ab_6__19_, ab_6__18_,
         ab_6__17_, ab_6__16_, ab_6__15_, ab_6__14_, ab_6__13_, ab_6__12_,
         ab_6__11_, ab_6__10_, ab_6__9_, ab_6__8_, ab_6__7_, ab_6__6_,
         ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_, ab_6__1_, ab_6__0_, ab_5__22_,
         ab_5__21_, ab_5__20_, ab_5__19_, ab_5__18_, ab_5__17_, ab_5__16_,
         ab_5__15_, ab_5__14_, ab_5__13_, ab_5__12_, ab_5__11_, ab_5__10_,
         ab_5__9_, ab_5__8_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__22_, ab_4__21_, ab_4__20_,
         ab_4__19_, ab_4__18_, ab_4__17_, ab_4__16_, ab_4__15_, ab_4__14_,
         ab_4__13_, ab_4__12_, ab_4__11_, ab_4__10_, ab_4__9_, ab_4__8_,
         ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_, ab_4__3_, ab_4__2_, ab_4__1_,
         ab_4__0_, ab_3__22_, ab_3__21_, ab_3__20_, ab_3__19_, ab_3__18_,
         ab_3__17_, ab_3__16_, ab_3__15_, ab_3__14_, ab_3__13_, ab_3__12_,
         ab_3__11_, ab_3__10_, ab_3__9_, ab_3__8_, ab_3__7_, ab_3__6_,
         ab_3__5_, ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__22_,
         ab_2__21_, ab_2__20_, ab_2__19_, ab_2__18_, ab_2__17_, ab_2__16_,
         ab_2__15_, ab_2__14_, ab_2__13_, ab_2__12_, ab_2__11_, ab_2__10_,
         ab_2__9_, ab_2__8_, ab_2__7_, ab_2__6_, ab_2__5_, ab_2__4_, ab_2__3_,
         ab_2__2_, ab_2__1_, ab_2__0_, ab_1__22_, ab_1__21_, ab_1__20_,
         ab_1__19_, ab_1__18_, ab_1__17_, ab_1__16_, ab_1__15_, ab_1__14_,
         ab_1__13_, ab_1__12_, ab_1__11_, ab_1__10_, ab_1__9_, ab_1__8_,
         ab_1__7_, ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_,
         ab_0__22_, ab_0__21_, ab_0__20_, ab_0__19_, ab_0__18_, ab_0__17_,
         ab_0__16_, ab_0__15_, ab_0__14_, ab_0__13_, ab_0__12_, ab_0__11_,
         ab_0__10_, ab_0__9_, ab_0__8_, ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_,
         ab_0__3_, ab_0__2_, CARRYB_23__22_, CARRYB_23__21_, CARRYB_23__20_,
         CARRYB_23__19_, CARRYB_23__18_, CARRYB_23__17_, CARRYB_23__16_,
         CARRYB_23__15_, CARRYB_23__14_, CARRYB_23__13_, CARRYB_23__12_,
         CARRYB_23__11_, CARRYB_23__10_, CARRYB_23__9_, CARRYB_23__8_,
         CARRYB_23__7_, CARRYB_23__6_, CARRYB_23__5_, CARRYB_23__4_,
         CARRYB_23__3_, CARRYB_23__2_, CARRYB_23__1_, CARRYB_23__0_,
         CARRYB_22__22_, CARRYB_22__21_, CARRYB_22__20_, CARRYB_22__19_,
         CARRYB_22__18_, CARRYB_22__17_, CARRYB_22__16_, CARRYB_22__15_,
         CARRYB_22__14_, CARRYB_22__13_, CARRYB_22__12_, CARRYB_22__11_,
         CARRYB_22__10_, CARRYB_22__9_, CARRYB_22__8_, CARRYB_22__7_,
         CARRYB_22__6_, CARRYB_22__5_, CARRYB_22__4_, CARRYB_22__3_,
         CARRYB_22__2_, CARRYB_22__1_, CARRYB_22__0_, CARRYB_21__22_,
         CARRYB_21__21_, CARRYB_21__20_, CARRYB_21__19_, CARRYB_21__18_,
         CARRYB_21__17_, CARRYB_21__16_, CARRYB_21__15_, CARRYB_21__14_,
         CARRYB_21__13_, CARRYB_21__12_, CARRYB_21__11_, CARRYB_21__10_,
         CARRYB_21__9_, CARRYB_21__8_, CARRYB_21__7_, CARRYB_21__6_,
         CARRYB_21__5_, CARRYB_21__4_, CARRYB_21__3_, CARRYB_21__2_,
         CARRYB_21__1_, CARRYB_21__0_, CARRYB_20__22_, CARRYB_20__21_,
         CARRYB_20__20_, CARRYB_20__19_, CARRYB_20__18_, CARRYB_20__17_,
         CARRYB_20__16_, CARRYB_20__15_, CARRYB_20__14_, CARRYB_20__13_,
         CARRYB_20__12_, CARRYB_20__11_, CARRYB_20__10_, CARRYB_20__9_,
         CARRYB_20__8_, CARRYB_20__7_, CARRYB_20__6_, CARRYB_20__5_,
         CARRYB_20__4_, CARRYB_20__3_, CARRYB_20__2_, CARRYB_20__1_,
         CARRYB_20__0_, CARRYB_19__22_, CARRYB_19__21_, CARRYB_19__20_,
         CARRYB_19__19_, CARRYB_19__18_, CARRYB_19__17_, CARRYB_19__16_,
         CARRYB_19__15_, CARRYB_19__14_, CARRYB_19__13_, CARRYB_19__12_,
         CARRYB_19__11_, CARRYB_19__10_, CARRYB_19__9_, CARRYB_19__8_,
         CARRYB_19__7_, CARRYB_19__6_, CARRYB_19__5_, CARRYB_19__4_,
         CARRYB_19__3_, CARRYB_19__2_, CARRYB_19__1_, CARRYB_19__0_,
         CARRYB_18__22_, CARRYB_18__21_, CARRYB_18__20_, CARRYB_18__19_,
         CARRYB_18__18_, CARRYB_18__17_, CARRYB_18__16_, CARRYB_18__15_,
         CARRYB_18__14_, CARRYB_18__13_, CARRYB_18__12_, CARRYB_18__11_,
         CARRYB_18__10_, CARRYB_18__9_, CARRYB_18__8_, CARRYB_18__7_,
         CARRYB_18__6_, CARRYB_18__5_, CARRYB_18__4_, CARRYB_18__3_,
         CARRYB_18__2_, CARRYB_18__1_, CARRYB_18__0_, CARRYB_17__22_,
         CARRYB_17__21_, CARRYB_17__20_, CARRYB_17__19_, CARRYB_17__18_,
         CARRYB_17__17_, CARRYB_17__16_, CARRYB_17__15_, CARRYB_17__14_,
         CARRYB_17__13_, CARRYB_17__12_, CARRYB_17__11_, CARRYB_17__10_,
         CARRYB_17__9_, CARRYB_17__8_, CARRYB_17__7_, CARRYB_17__6_,
         CARRYB_17__5_, CARRYB_17__4_, CARRYB_17__3_, CARRYB_17__2_,
         CARRYB_17__1_, CARRYB_17__0_, CARRYB_16__22_, CARRYB_16__21_,
         CARRYB_16__20_, CARRYB_16__19_, CARRYB_16__18_, CARRYB_16__17_,
         CARRYB_16__16_, CARRYB_16__15_, CARRYB_16__14_, CARRYB_16__13_,
         CARRYB_16__12_, CARRYB_16__11_, CARRYB_16__10_, CARRYB_16__9_,
         CARRYB_16__8_, CARRYB_16__7_, CARRYB_16__6_, CARRYB_16__5_,
         CARRYB_16__4_, CARRYB_16__3_, CARRYB_16__2_, CARRYB_16__1_,
         CARRYB_16__0_, CARRYB_15__22_, CARRYB_15__21_, CARRYB_15__20_,
         CARRYB_15__19_, CARRYB_15__18_, CARRYB_15__17_, CARRYB_15__16_,
         CARRYB_15__15_, CARRYB_15__14_, CARRYB_15__13_, CARRYB_15__12_,
         CARRYB_15__11_, CARRYB_15__10_, CARRYB_15__9_, CARRYB_15__8_,
         CARRYB_15__7_, CARRYB_15__6_, CARRYB_15__5_, CARRYB_15__4_,
         CARRYB_15__3_, CARRYB_15__2_, CARRYB_15__1_, CARRYB_15__0_,
         CARRYB_14__22_, CARRYB_14__21_, CARRYB_14__20_, CARRYB_14__19_,
         CARRYB_14__18_, CARRYB_14__17_, CARRYB_14__16_, CARRYB_14__15_,
         CARRYB_14__14_, CARRYB_14__13_, CARRYB_14__12_, CARRYB_14__11_,
         CARRYB_14__10_, CARRYB_14__9_, CARRYB_14__8_, CARRYB_14__7_,
         CARRYB_14__6_, CARRYB_14__5_, CARRYB_14__4_, CARRYB_14__3_,
         CARRYB_14__2_, CARRYB_14__1_, CARRYB_14__0_, CARRYB_13__22_,
         CARRYB_13__21_, CARRYB_13__20_, CARRYB_13__19_, CARRYB_13__18_,
         CARRYB_13__17_, CARRYB_13__16_, CARRYB_13__15_, CARRYB_13__14_,
         CARRYB_13__13_, CARRYB_13__12_, CARRYB_13__11_, CARRYB_13__10_,
         CARRYB_13__9_, CARRYB_13__8_, CARRYB_13__7_, CARRYB_13__6_,
         CARRYB_13__5_, CARRYB_13__4_, CARRYB_13__3_, CARRYB_13__2_,
         CARRYB_13__1_, CARRYB_13__0_, CARRYB_12__22_, CARRYB_12__21_,
         CARRYB_12__20_, CARRYB_12__19_, CARRYB_12__18_, CARRYB_12__17_,
         CARRYB_12__16_, CARRYB_12__15_, CARRYB_12__14_, CARRYB_12__13_,
         CARRYB_12__12_, CARRYB_12__11_, CARRYB_12__10_, CARRYB_12__9_,
         CARRYB_12__8_, CARRYB_12__7_, CARRYB_12__6_, CARRYB_12__5_,
         CARRYB_12__4_, CARRYB_12__3_, CARRYB_12__2_, CARRYB_12__1_,
         CARRYB_12__0_, CARRYB_11__22_, CARRYB_11__21_, CARRYB_11__20_,
         CARRYB_11__19_, CARRYB_11__18_, CARRYB_11__17_, CARRYB_11__16_,
         CARRYB_11__15_, CARRYB_11__14_, CARRYB_11__13_, CARRYB_11__12_,
         CARRYB_11__11_, CARRYB_11__10_, CARRYB_11__9_, CARRYB_11__8_,
         CARRYB_11__7_, CARRYB_11__6_, CARRYB_11__5_, CARRYB_11__4_,
         CARRYB_11__3_, CARRYB_11__2_, CARRYB_11__1_, CARRYB_11__0_,
         CARRYB_10__22_, CARRYB_10__21_, CARRYB_10__20_, CARRYB_10__19_,
         CARRYB_10__18_, CARRYB_10__17_, CARRYB_10__16_, CARRYB_10__15_,
         CARRYB_10__14_, CARRYB_10__13_, CARRYB_10__12_, CARRYB_10__11_,
         CARRYB_10__10_, CARRYB_10__9_, CARRYB_10__8_, CARRYB_10__7_,
         CARRYB_10__6_, CARRYB_10__5_, CARRYB_10__4_, CARRYB_10__3_,
         CARRYB_10__2_, CARRYB_10__1_, CARRYB_10__0_, CARRYB_9__22_,
         CARRYB_9__21_, CARRYB_9__20_, CARRYB_9__19_, CARRYB_9__18_,
         CARRYB_9__17_, CARRYB_9__16_, CARRYB_9__15_, CARRYB_9__14_,
         CARRYB_9__13_, CARRYB_9__12_, CARRYB_9__11_, CARRYB_9__10_,
         CARRYB_9__9_, CARRYB_9__8_, CARRYB_9__7_, CARRYB_9__6_, CARRYB_9__5_,
         CARRYB_9__4_, CARRYB_9__3_, CARRYB_9__2_, CARRYB_9__1_, CARRYB_9__0_,
         CARRYB_8__22_, CARRYB_8__21_, CARRYB_8__20_, CARRYB_8__19_,
         CARRYB_8__18_, CARRYB_8__17_, CARRYB_8__16_, CARRYB_8__15_,
         CARRYB_8__14_, CARRYB_8__13_, CARRYB_8__12_, CARRYB_8__11_,
         CARRYB_8__10_, CARRYB_8__9_, CARRYB_8__8_, CARRYB_8__7_, CARRYB_8__6_,
         CARRYB_8__5_, CARRYB_8__4_, CARRYB_8__3_, CARRYB_8__2_, CARRYB_8__1_,
         CARRYB_8__0_, CARRYB_7__22_, CARRYB_7__21_, CARRYB_7__20_,
         CARRYB_7__19_, CARRYB_7__18_, CARRYB_7__17_, CARRYB_7__16_,
         CARRYB_7__15_, CARRYB_7__14_, CARRYB_7__13_, CARRYB_7__12_,
         CARRYB_7__11_, CARRYB_7__10_, CARRYB_7__9_, CARRYB_7__8_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__22_,
         CARRYB_6__21_, CARRYB_6__20_, CARRYB_6__19_, CARRYB_6__18_,
         CARRYB_6__17_, CARRYB_6__16_, CARRYB_6__15_, CARRYB_6__14_,
         CARRYB_6__13_, CARRYB_6__12_, CARRYB_6__11_, CARRYB_6__10_,
         CARRYB_6__9_, CARRYB_6__8_, CARRYB_6__7_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__22_, CARRYB_5__21_, CARRYB_5__20_, CARRYB_5__19_,
         CARRYB_5__18_, CARRYB_5__17_, CARRYB_5__16_, CARRYB_5__15_,
         CARRYB_5__14_, CARRYB_5__13_, CARRYB_5__12_, CARRYB_5__11_,
         CARRYB_5__10_, CARRYB_5__9_, CARRYB_5__8_, CARRYB_5__7_, CARRYB_5__6_,
         CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_, CARRYB_5__1_,
         CARRYB_5__0_, CARRYB_4__22_, CARRYB_4__21_, CARRYB_4__20_,
         CARRYB_4__19_, CARRYB_4__18_, CARRYB_4__17_, CARRYB_4__16_,
         CARRYB_4__15_, CARRYB_4__14_, CARRYB_4__13_, CARRYB_4__12_,
         CARRYB_4__11_, CARRYB_4__10_, CARRYB_4__9_, CARRYB_4__8_,
         CARRYB_4__7_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_, CARRYB_4__3_,
         CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__22_,
         CARRYB_3__21_, CARRYB_3__20_, CARRYB_3__19_, CARRYB_3__18_,
         CARRYB_3__17_, CARRYB_3__16_, CARRYB_3__15_, CARRYB_3__14_,
         CARRYB_3__13_, CARRYB_3__12_, CARRYB_3__11_, CARRYB_3__10_,
         CARRYB_3__9_, CARRYB_3__8_, CARRYB_3__7_, CARRYB_3__6_, CARRYB_3__5_,
         CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_, CARRYB_3__0_,
         CARRYB_2__22_, CARRYB_2__21_, CARRYB_2__20_, CARRYB_2__19_,
         CARRYB_2__18_, CARRYB_2__17_, CARRYB_2__16_, CARRYB_2__15_,
         CARRYB_2__14_, CARRYB_2__13_, CARRYB_2__12_, CARRYB_2__11_,
         CARRYB_2__10_, CARRYB_2__9_, CARRYB_2__8_, CARRYB_2__7_, CARRYB_2__6_,
         CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_, CARRYB_2__2_, CARRYB_2__1_,
         CARRYB_2__0_, CARRYB_1__0_, SUMB_23__22_, SUMB_23__21_, SUMB_23__20_,
         SUMB_23__19_, SUMB_23__18_, SUMB_23__17_, SUMB_23__16_, SUMB_23__15_,
         SUMB_23__14_, SUMB_23__13_, SUMB_23__12_, SUMB_23__11_, SUMB_23__10_,
         SUMB_23__9_, SUMB_23__8_, SUMB_23__7_, SUMB_23__6_, SUMB_23__5_,
         SUMB_23__4_, SUMB_23__3_, SUMB_23__2_, SUMB_23__1_, SUMB_23__0_,
         SUMB_22__22_, SUMB_22__21_, SUMB_22__20_, SUMB_22__19_, SUMB_22__18_,
         SUMB_22__17_, SUMB_22__16_, SUMB_22__15_, SUMB_22__14_, SUMB_22__13_,
         SUMB_22__12_, SUMB_22__11_, SUMB_22__10_, SUMB_22__9_, SUMB_22__8_,
         SUMB_22__7_, SUMB_22__6_, SUMB_22__5_, SUMB_22__4_, SUMB_22__3_,
         SUMB_22__2_, SUMB_22__1_, SUMB_21__22_, SUMB_21__21_, SUMB_21__20_,
         SUMB_21__19_, SUMB_21__18_, SUMB_21__17_, SUMB_21__16_, SUMB_21__15_,
         SUMB_21__14_, SUMB_21__13_, SUMB_21__12_, SUMB_21__11_, SUMB_21__10_,
         SUMB_21__9_, SUMB_21__8_, SUMB_21__7_, SUMB_21__6_, SUMB_21__5_,
         SUMB_21__4_, SUMB_21__3_, SUMB_21__2_, SUMB_21__1_, SUMB_20__22_,
         SUMB_20__21_, SUMB_20__20_, SUMB_20__19_, SUMB_20__18_, SUMB_20__17_,
         SUMB_20__16_, SUMB_20__15_, SUMB_20__14_, SUMB_20__13_, SUMB_20__12_,
         SUMB_20__11_, SUMB_20__10_, SUMB_20__9_, SUMB_20__8_, SUMB_20__7_,
         SUMB_20__6_, SUMB_20__5_, SUMB_20__4_, SUMB_20__3_, SUMB_20__2_,
         SUMB_20__1_, SUMB_19__22_, SUMB_19__21_, SUMB_19__20_, SUMB_19__19_,
         SUMB_19__18_, SUMB_19__17_, SUMB_19__16_, SUMB_19__15_, SUMB_19__14_,
         SUMB_19__13_, SUMB_19__12_, SUMB_19__11_, SUMB_19__10_, SUMB_19__9_,
         SUMB_19__8_, SUMB_19__7_, SUMB_19__6_, SUMB_19__5_, SUMB_19__4_,
         SUMB_19__3_, SUMB_19__2_, SUMB_19__1_, SUMB_18__22_, SUMB_18__21_,
         SUMB_18__20_, SUMB_18__19_, SUMB_18__18_, SUMB_18__17_, SUMB_18__16_,
         SUMB_18__15_, SUMB_18__14_, SUMB_18__13_, SUMB_18__12_, SUMB_18__11_,
         SUMB_18__10_, SUMB_18__9_, SUMB_18__8_, SUMB_18__7_, SUMB_18__6_,
         SUMB_18__5_, SUMB_18__4_, SUMB_18__3_, SUMB_18__2_, SUMB_18__1_,
         SUMB_17__22_, SUMB_17__21_, SUMB_17__20_, SUMB_17__19_, SUMB_17__18_,
         SUMB_17__17_, SUMB_17__16_, SUMB_17__15_, SUMB_17__14_, SUMB_17__13_,
         SUMB_17__12_, SUMB_17__11_, SUMB_17__10_, SUMB_17__9_, SUMB_17__8_,
         SUMB_17__7_, SUMB_17__6_, SUMB_17__5_, SUMB_17__4_, SUMB_17__3_,
         SUMB_17__2_, SUMB_17__1_, SUMB_16__22_, SUMB_16__21_, SUMB_16__20_,
         SUMB_16__19_, SUMB_16__18_, SUMB_16__17_, SUMB_16__16_, SUMB_16__15_,
         SUMB_16__14_, SUMB_16__13_, SUMB_16__12_, SUMB_16__11_, SUMB_16__10_,
         SUMB_16__9_, SUMB_16__8_, SUMB_16__7_, SUMB_16__6_, SUMB_16__5_,
         SUMB_16__4_, SUMB_16__3_, SUMB_16__2_, SUMB_16__1_, SUMB_15__22_,
         SUMB_15__21_, SUMB_15__20_, SUMB_15__19_, SUMB_15__18_, SUMB_15__17_,
         SUMB_15__16_, SUMB_15__15_, SUMB_15__14_, SUMB_15__13_, SUMB_15__12_,
         SUMB_15__11_, SUMB_15__10_, SUMB_15__9_, SUMB_15__8_, SUMB_15__7_,
         SUMB_15__6_, SUMB_15__5_, SUMB_15__4_, SUMB_15__3_, SUMB_15__2_,
         SUMB_15__1_, SUMB_14__22_, SUMB_14__21_, SUMB_14__20_, SUMB_14__19_,
         SUMB_14__18_, SUMB_14__17_, SUMB_14__16_, SUMB_14__15_, SUMB_14__14_,
         SUMB_14__13_, SUMB_14__12_, SUMB_14__11_, SUMB_14__10_, SUMB_14__9_,
         SUMB_14__8_, SUMB_14__7_, SUMB_14__6_, SUMB_14__5_, SUMB_14__4_,
         SUMB_14__3_, SUMB_14__2_, SUMB_14__1_, SUMB_13__22_, SUMB_13__21_,
         SUMB_13__20_, SUMB_13__19_, SUMB_13__18_, SUMB_13__17_, SUMB_13__16_,
         SUMB_13__15_, SUMB_13__14_, SUMB_13__13_, SUMB_13__12_, SUMB_13__11_,
         SUMB_13__10_, SUMB_13__9_, SUMB_13__8_, SUMB_13__7_, SUMB_13__6_,
         SUMB_13__5_, SUMB_13__4_, SUMB_13__3_, SUMB_13__2_, SUMB_13__1_,
         SUMB_12__22_, SUMB_12__21_, SUMB_12__20_, SUMB_12__19_, SUMB_12__18_,
         SUMB_12__17_, SUMB_12__16_, SUMB_12__15_, SUMB_12__14_, SUMB_12__13_,
         SUMB_12__12_, SUMB_12__11_, SUMB_12__10_, SUMB_12__9_, SUMB_12__8_,
         SUMB_12__7_, SUMB_12__6_, SUMB_12__5_, SUMB_12__4_, SUMB_12__3_,
         SUMB_12__2_, SUMB_12__1_, SUMB_11__22_, SUMB_11__21_, SUMB_11__20_,
         SUMB_11__19_, SUMB_11__18_, SUMB_11__17_, SUMB_11__16_, SUMB_11__15_,
         SUMB_11__14_, SUMB_11__13_, SUMB_11__12_, SUMB_11__11_, SUMB_11__10_,
         SUMB_11__9_, SUMB_11__8_, SUMB_11__7_, SUMB_11__6_, SUMB_11__5_,
         SUMB_11__4_, SUMB_11__3_, SUMB_11__2_, SUMB_11__1_, SUMB_10__22_,
         SUMB_10__21_, SUMB_10__20_, SUMB_10__19_, SUMB_10__18_, SUMB_10__17_,
         SUMB_10__16_, SUMB_10__15_, SUMB_10__14_, SUMB_10__13_, SUMB_10__12_,
         SUMB_10__11_, SUMB_10__10_, SUMB_10__9_, SUMB_10__8_, SUMB_10__7_,
         SUMB_10__6_, SUMB_10__5_, SUMB_10__4_, SUMB_10__3_, SUMB_10__2_,
         SUMB_10__1_, SUMB_9__22_, SUMB_9__21_, SUMB_9__20_, SUMB_9__19_,
         SUMB_9__18_, SUMB_9__17_, SUMB_9__16_, SUMB_9__15_, SUMB_9__14_,
         SUMB_9__13_, SUMB_9__12_, SUMB_9__11_, SUMB_9__10_, SUMB_9__9_,
         SUMB_9__8_, SUMB_9__7_, SUMB_9__6_, SUMB_9__5_, SUMB_9__4_,
         SUMB_9__3_, SUMB_9__2_, SUMB_9__1_, SUMB_8__22_, SUMB_8__21_,
         SUMB_8__20_, SUMB_8__19_, SUMB_8__18_, SUMB_8__17_, SUMB_8__16_,
         SUMB_8__15_, SUMB_8__14_, SUMB_8__13_, SUMB_8__12_, SUMB_8__11_,
         SUMB_8__10_, SUMB_8__9_, SUMB_8__8_, SUMB_8__7_, SUMB_8__6_,
         SUMB_8__5_, SUMB_8__4_, SUMB_8__3_, SUMB_8__2_, SUMB_8__1_,
         SUMB_7__22_, SUMB_7__21_, SUMB_7__20_, SUMB_7__19_, SUMB_7__18_,
         SUMB_7__17_, SUMB_7__16_, SUMB_7__15_, SUMB_7__14_, SUMB_7__13_,
         SUMB_7__12_, SUMB_7__11_, SUMB_7__10_, SUMB_7__9_, SUMB_7__8_,
         SUMB_7__7_, SUMB_7__6_, SUMB_7__5_, SUMB_7__4_, SUMB_7__3_,
         SUMB_7__2_, SUMB_7__1_, SUMB_6__22_, SUMB_6__21_, SUMB_6__20_,
         SUMB_6__19_, SUMB_6__18_, SUMB_6__17_, SUMB_6__16_, SUMB_6__15_,
         SUMB_6__14_, SUMB_6__13_, SUMB_6__12_, SUMB_6__11_, SUMB_6__10_,
         SUMB_6__9_, SUMB_6__8_, SUMB_6__7_, SUMB_6__6_, SUMB_6__5_,
         SUMB_6__4_, SUMB_6__3_, SUMB_6__2_, SUMB_6__1_, SUMB_5__22_,
         SUMB_5__21_, SUMB_5__20_, SUMB_5__19_, SUMB_5__18_, SUMB_5__17_,
         SUMB_5__16_, SUMB_5__15_, SUMB_5__14_, SUMB_5__13_, SUMB_5__12_,
         SUMB_5__11_, SUMB_5__10_, SUMB_5__9_, SUMB_5__8_, SUMB_5__7_,
         SUMB_5__6_, SUMB_5__5_, SUMB_5__4_, SUMB_5__3_, SUMB_5__2_,
         SUMB_5__1_, SUMB_4__22_, SUMB_4__21_, SUMB_4__20_, SUMB_4__19_,
         SUMB_4__18_, SUMB_4__17_, SUMB_4__16_, SUMB_4__15_, SUMB_4__14_,
         SUMB_4__13_, SUMB_4__12_, SUMB_4__11_, SUMB_4__10_, SUMB_4__9_,
         SUMB_4__8_, SUMB_4__7_, SUMB_4__6_, SUMB_4__5_, SUMB_4__4_,
         SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__22_, SUMB_3__21_,
         SUMB_3__20_, SUMB_3__19_, SUMB_3__18_, SUMB_3__17_, SUMB_3__16_,
         SUMB_3__15_, SUMB_3__14_, SUMB_3__13_, SUMB_3__12_, SUMB_3__11_,
         SUMB_3__10_, SUMB_3__9_, SUMB_3__8_, SUMB_3__7_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__22_, SUMB_2__21_, SUMB_2__20_, SUMB_2__19_, SUMB_2__18_,
         SUMB_2__17_, SUMB_2__16_, SUMB_2__15_, SUMB_2__14_, SUMB_2__13_,
         SUMB_2__12_, SUMB_2__11_, SUMB_2__10_, SUMB_2__9_, SUMB_2__8_,
         SUMB_2__7_, SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_,
         SUMB_2__2_, SUMB_2__1_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_,
         A1_15_, A1_14_, A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_,
         A1_6_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7,
         SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9,
         SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11,
         SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13,
         SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15,
         SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17,
         SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19,
         SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21;

  FA_X1 S4_0 ( .A(B[0]), .B(CARRYB_22__0_), .CI(SUMB_22__1_), .CO(
        CARRYB_23__0_), .S(SUMB_23__0_) );
  FA_X1 S4_1 ( .A(B[1]), .B(CARRYB_22__1_), .CI(SUMB_22__2_), .CO(
        CARRYB_23__1_), .S(SUMB_23__1_) );
  FA_X1 S4_2 ( .A(B[2]), .B(CARRYB_22__2_), .CI(SUMB_22__3_), .CO(
        CARRYB_23__2_), .S(SUMB_23__2_) );
  FA_X1 S4_3 ( .A(B[3]), .B(CARRYB_22__3_), .CI(SUMB_22__4_), .CO(
        CARRYB_23__3_), .S(SUMB_23__3_) );
  FA_X1 S4_4 ( .A(B[4]), .B(CARRYB_22__4_), .CI(SUMB_22__5_), .CO(
        CARRYB_23__4_), .S(SUMB_23__4_) );
  FA_X1 S4_5 ( .A(B[5]), .B(CARRYB_22__5_), .CI(SUMB_22__6_), .CO(
        CARRYB_23__5_), .S(SUMB_23__5_) );
  FA_X1 S4_6 ( .A(B[6]), .B(CARRYB_22__6_), .CI(SUMB_22__7_), .CO(
        CARRYB_23__6_), .S(SUMB_23__6_) );
  FA_X1 S4_7 ( .A(B[7]), .B(CARRYB_22__7_), .CI(SUMB_22__8_), .CO(
        CARRYB_23__7_), .S(SUMB_23__7_) );
  FA_X1 S4_8 ( .A(B[8]), .B(CARRYB_22__8_), .CI(SUMB_22__9_), .CO(
        CARRYB_23__8_), .S(SUMB_23__8_) );
  FA_X1 S4_9 ( .A(B[9]), .B(CARRYB_22__9_), .CI(SUMB_22__10_), .CO(
        CARRYB_23__9_), .S(SUMB_23__9_) );
  FA_X1 S4_10 ( .A(B[10]), .B(CARRYB_22__10_), .CI(SUMB_22__11_), .CO(
        CARRYB_23__10_), .S(SUMB_23__10_) );
  FA_X1 S4_11 ( .A(B[11]), .B(CARRYB_22__11_), .CI(SUMB_22__12_), .CO(
        CARRYB_23__11_), .S(SUMB_23__11_) );
  FA_X1 S4_12 ( .A(B[12]), .B(CARRYB_22__12_), .CI(SUMB_22__13_), .CO(
        CARRYB_23__12_), .S(SUMB_23__12_) );
  FA_X1 S4_13 ( .A(B[13]), .B(CARRYB_22__13_), .CI(SUMB_22__14_), .CO(
        CARRYB_23__13_), .S(SUMB_23__13_) );
  FA_X1 S4_14 ( .A(B[14]), .B(CARRYB_22__14_), .CI(SUMB_22__15_), .CO(
        CARRYB_23__14_), .S(SUMB_23__14_) );
  FA_X1 S4_15 ( .A(B[15]), .B(CARRYB_22__15_), .CI(SUMB_22__16_), .CO(
        CARRYB_23__15_), .S(SUMB_23__15_) );
  FA_X1 S4_16 ( .A(B[16]), .B(CARRYB_22__16_), .CI(SUMB_22__17_), .CO(
        CARRYB_23__16_), .S(SUMB_23__16_) );
  FA_X1 S4_17 ( .A(B[17]), .B(CARRYB_22__17_), .CI(SUMB_22__18_), .CO(
        CARRYB_23__17_), .S(SUMB_23__17_) );
  FA_X1 S4_18 ( .A(B[18]), .B(CARRYB_22__18_), .CI(SUMB_22__19_), .CO(
        CARRYB_23__18_), .S(SUMB_23__18_) );
  FA_X1 S4_19 ( .A(B[19]), .B(CARRYB_22__19_), .CI(SUMB_22__20_), .CO(
        CARRYB_23__19_), .S(SUMB_23__19_) );
  FA_X1 S4_20 ( .A(B[20]), .B(CARRYB_22__20_), .CI(SUMB_22__21_), .CO(
        CARRYB_23__20_), .S(SUMB_23__20_) );
  FA_X1 S4_21 ( .A(B[21]), .B(CARRYB_22__21_), .CI(SUMB_22__22_), .CO(
        CARRYB_23__21_), .S(SUMB_23__21_) );
  FA_X1 S5_22 ( .A(B[22]), .B(CARRYB_22__22_), .CI(A[22]), .CO(CARRYB_23__22_), 
        .S(SUMB_23__22_) );
  FA_X1 S1_22_0 ( .A(ab_22__0_), .B(CARRYB_21__0_), .CI(SUMB_21__1_), .CO(
        CARRYB_22__0_), .S(A1_20_) );
  FA_X1 S2_22_1 ( .A(ab_22__1_), .B(CARRYB_21__1_), .CI(SUMB_21__2_), .CO(
        CARRYB_22__1_), .S(SUMB_22__1_) );
  FA_X1 S2_22_2 ( .A(ab_22__2_), .B(CARRYB_21__2_), .CI(SUMB_21__3_), .CO(
        CARRYB_22__2_), .S(SUMB_22__2_) );
  FA_X1 S2_22_3 ( .A(ab_22__3_), .B(CARRYB_21__3_), .CI(SUMB_21__4_), .CO(
        CARRYB_22__3_), .S(SUMB_22__3_) );
  FA_X1 S2_22_4 ( .A(ab_22__4_), .B(CARRYB_21__4_), .CI(SUMB_21__5_), .CO(
        CARRYB_22__4_), .S(SUMB_22__4_) );
  FA_X1 S2_22_5 ( .A(ab_22__5_), .B(CARRYB_21__5_), .CI(SUMB_21__6_), .CO(
        CARRYB_22__5_), .S(SUMB_22__5_) );
  FA_X1 S2_22_6 ( .A(ab_22__6_), .B(CARRYB_21__6_), .CI(SUMB_21__7_), .CO(
        CARRYB_22__6_), .S(SUMB_22__6_) );
  FA_X1 S2_22_7 ( .A(ab_22__7_), .B(CARRYB_21__7_), .CI(SUMB_21__8_), .CO(
        CARRYB_22__7_), .S(SUMB_22__7_) );
  FA_X1 S2_22_8 ( .A(ab_22__8_), .B(CARRYB_21__8_), .CI(SUMB_21__9_), .CO(
        CARRYB_22__8_), .S(SUMB_22__8_) );
  FA_X1 S2_22_9 ( .A(ab_22__9_), .B(CARRYB_21__9_), .CI(SUMB_21__10_), .CO(
        CARRYB_22__9_), .S(SUMB_22__9_) );
  FA_X1 S2_22_10 ( .A(ab_22__10_), .B(CARRYB_21__10_), .CI(SUMB_21__11_), .CO(
        CARRYB_22__10_), .S(SUMB_22__10_) );
  FA_X1 S2_22_11 ( .A(ab_22__11_), .B(CARRYB_21__11_), .CI(SUMB_21__12_), .CO(
        CARRYB_22__11_), .S(SUMB_22__11_) );
  FA_X1 S2_22_12 ( .A(ab_22__12_), .B(CARRYB_21__12_), .CI(SUMB_21__13_), .CO(
        CARRYB_22__12_), .S(SUMB_22__12_) );
  FA_X1 S2_22_13 ( .A(ab_22__13_), .B(CARRYB_21__13_), .CI(SUMB_21__14_), .CO(
        CARRYB_22__13_), .S(SUMB_22__13_) );
  FA_X1 S2_22_14 ( .A(ab_22__14_), .B(CARRYB_21__14_), .CI(SUMB_21__15_), .CO(
        CARRYB_22__14_), .S(SUMB_22__14_) );
  FA_X1 S2_22_15 ( .A(ab_22__15_), .B(CARRYB_21__15_), .CI(SUMB_21__16_), .CO(
        CARRYB_22__15_), .S(SUMB_22__15_) );
  FA_X1 S2_22_16 ( .A(ab_22__16_), .B(CARRYB_21__16_), .CI(SUMB_21__17_), .CO(
        CARRYB_22__16_), .S(SUMB_22__16_) );
  FA_X1 S2_22_17 ( .A(ab_22__17_), .B(CARRYB_21__17_), .CI(SUMB_21__18_), .CO(
        CARRYB_22__17_), .S(SUMB_22__17_) );
  FA_X1 S2_22_18 ( .A(ab_22__18_), .B(CARRYB_21__18_), .CI(SUMB_21__19_), .CO(
        CARRYB_22__18_), .S(SUMB_22__18_) );
  FA_X1 S2_22_19 ( .A(ab_22__19_), .B(CARRYB_21__19_), .CI(SUMB_21__20_), .CO(
        CARRYB_22__19_), .S(SUMB_22__19_) );
  FA_X1 S2_22_20 ( .A(ab_22__20_), .B(CARRYB_21__20_), .CI(SUMB_21__21_), .CO(
        CARRYB_22__20_), .S(SUMB_22__20_) );
  FA_X1 S2_22_21 ( .A(ab_22__21_), .B(CARRYB_21__21_), .CI(SUMB_21__22_), .CO(
        CARRYB_22__21_), .S(SUMB_22__21_) );
  FA_X1 S3_22_22 ( .A(ab_22__22_), .B(CARRYB_21__22_), .CI(A[21]), .CO(
        CARRYB_22__22_), .S(SUMB_22__22_) );
  FA_X1 S1_21_0 ( .A(ab_21__0_), .B(CARRYB_20__0_), .CI(SUMB_20__1_), .CO(
        CARRYB_21__0_), .S(A1_19_) );
  FA_X1 S2_21_1 ( .A(ab_21__1_), .B(CARRYB_20__1_), .CI(SUMB_20__2_), .CO(
        CARRYB_21__1_), .S(SUMB_21__1_) );
  FA_X1 S2_21_2 ( .A(ab_21__2_), .B(CARRYB_20__2_), .CI(SUMB_20__3_), .CO(
        CARRYB_21__2_), .S(SUMB_21__2_) );
  FA_X1 S2_21_3 ( .A(ab_21__3_), .B(CARRYB_20__3_), .CI(SUMB_20__4_), .CO(
        CARRYB_21__3_), .S(SUMB_21__3_) );
  FA_X1 S2_21_4 ( .A(ab_21__4_), .B(CARRYB_20__4_), .CI(SUMB_20__5_), .CO(
        CARRYB_21__4_), .S(SUMB_21__4_) );
  FA_X1 S2_21_5 ( .A(ab_21__5_), .B(CARRYB_20__5_), .CI(SUMB_20__6_), .CO(
        CARRYB_21__5_), .S(SUMB_21__5_) );
  FA_X1 S2_21_6 ( .A(ab_21__6_), .B(CARRYB_20__6_), .CI(SUMB_20__7_), .CO(
        CARRYB_21__6_), .S(SUMB_21__6_) );
  FA_X1 S2_21_7 ( .A(ab_21__7_), .B(CARRYB_20__7_), .CI(SUMB_20__8_), .CO(
        CARRYB_21__7_), .S(SUMB_21__7_) );
  FA_X1 S2_21_8 ( .A(ab_21__8_), .B(CARRYB_20__8_), .CI(SUMB_20__9_), .CO(
        CARRYB_21__8_), .S(SUMB_21__8_) );
  FA_X1 S2_21_9 ( .A(ab_21__9_), .B(CARRYB_20__9_), .CI(SUMB_20__10_), .CO(
        CARRYB_21__9_), .S(SUMB_21__9_) );
  FA_X1 S2_21_10 ( .A(ab_21__10_), .B(CARRYB_20__10_), .CI(SUMB_20__11_), .CO(
        CARRYB_21__10_), .S(SUMB_21__10_) );
  FA_X1 S2_21_11 ( .A(ab_21__11_), .B(CARRYB_20__11_), .CI(SUMB_20__12_), .CO(
        CARRYB_21__11_), .S(SUMB_21__11_) );
  FA_X1 S2_21_12 ( .A(ab_21__12_), .B(CARRYB_20__12_), .CI(SUMB_20__13_), .CO(
        CARRYB_21__12_), .S(SUMB_21__12_) );
  FA_X1 S2_21_13 ( .A(ab_21__13_), .B(CARRYB_20__13_), .CI(SUMB_20__14_), .CO(
        CARRYB_21__13_), .S(SUMB_21__13_) );
  FA_X1 S2_21_14 ( .A(ab_21__14_), .B(CARRYB_20__14_), .CI(SUMB_20__15_), .CO(
        CARRYB_21__14_), .S(SUMB_21__14_) );
  FA_X1 S2_21_15 ( .A(ab_21__15_), .B(CARRYB_20__15_), .CI(SUMB_20__16_), .CO(
        CARRYB_21__15_), .S(SUMB_21__15_) );
  FA_X1 S2_21_16 ( .A(ab_21__16_), .B(CARRYB_20__16_), .CI(SUMB_20__17_), .CO(
        CARRYB_21__16_), .S(SUMB_21__16_) );
  FA_X1 S2_21_17 ( .A(ab_21__17_), .B(CARRYB_20__17_), .CI(SUMB_20__18_), .CO(
        CARRYB_21__17_), .S(SUMB_21__17_) );
  FA_X1 S2_21_18 ( .A(ab_21__18_), .B(CARRYB_20__18_), .CI(SUMB_20__19_), .CO(
        CARRYB_21__18_), .S(SUMB_21__18_) );
  FA_X1 S2_21_19 ( .A(ab_21__19_), .B(CARRYB_20__19_), .CI(SUMB_20__20_), .CO(
        CARRYB_21__19_), .S(SUMB_21__19_) );
  FA_X1 S2_21_20 ( .A(ab_21__20_), .B(CARRYB_20__20_), .CI(SUMB_20__21_), .CO(
        CARRYB_21__20_), .S(SUMB_21__20_) );
  FA_X1 S2_21_21 ( .A(ab_21__21_), .B(CARRYB_20__21_), .CI(SUMB_20__22_), .CO(
        CARRYB_21__21_), .S(SUMB_21__21_) );
  FA_X1 S3_21_22 ( .A(ab_21__22_), .B(CARRYB_20__22_), .CI(A[20]), .CO(
        CARRYB_21__22_), .S(SUMB_21__22_) );
  FA_X1 S1_20_0 ( .A(ab_20__0_), .B(CARRYB_19__0_), .CI(SUMB_19__1_), .CO(
        CARRYB_20__0_), .S(A1_18_) );
  FA_X1 S2_20_1 ( .A(ab_20__1_), .B(CARRYB_19__1_), .CI(SUMB_19__2_), .CO(
        CARRYB_20__1_), .S(SUMB_20__1_) );
  FA_X1 S2_20_2 ( .A(ab_20__2_), .B(CARRYB_19__2_), .CI(SUMB_19__3_), .CO(
        CARRYB_20__2_), .S(SUMB_20__2_) );
  FA_X1 S2_20_3 ( .A(ab_20__3_), .B(CARRYB_19__3_), .CI(SUMB_19__4_), .CO(
        CARRYB_20__3_), .S(SUMB_20__3_) );
  FA_X1 S2_20_4 ( .A(ab_20__4_), .B(CARRYB_19__4_), .CI(SUMB_19__5_), .CO(
        CARRYB_20__4_), .S(SUMB_20__4_) );
  FA_X1 S2_20_5 ( .A(ab_20__5_), .B(CARRYB_19__5_), .CI(SUMB_19__6_), .CO(
        CARRYB_20__5_), .S(SUMB_20__5_) );
  FA_X1 S2_20_6 ( .A(ab_20__6_), .B(CARRYB_19__6_), .CI(SUMB_19__7_), .CO(
        CARRYB_20__6_), .S(SUMB_20__6_) );
  FA_X1 S2_20_7 ( .A(ab_20__7_), .B(CARRYB_19__7_), .CI(SUMB_19__8_), .CO(
        CARRYB_20__7_), .S(SUMB_20__7_) );
  FA_X1 S2_20_8 ( .A(ab_20__8_), .B(CARRYB_19__8_), .CI(SUMB_19__9_), .CO(
        CARRYB_20__8_), .S(SUMB_20__8_) );
  FA_X1 S2_20_9 ( .A(ab_20__9_), .B(CARRYB_19__9_), .CI(SUMB_19__10_), .CO(
        CARRYB_20__9_), .S(SUMB_20__9_) );
  FA_X1 S2_20_10 ( .A(ab_20__10_), .B(CARRYB_19__10_), .CI(SUMB_19__11_), .CO(
        CARRYB_20__10_), .S(SUMB_20__10_) );
  FA_X1 S2_20_11 ( .A(ab_20__11_), .B(CARRYB_19__11_), .CI(SUMB_19__12_), .CO(
        CARRYB_20__11_), .S(SUMB_20__11_) );
  FA_X1 S2_20_12 ( .A(ab_20__12_), .B(CARRYB_19__12_), .CI(SUMB_19__13_), .CO(
        CARRYB_20__12_), .S(SUMB_20__12_) );
  FA_X1 S2_20_13 ( .A(ab_20__13_), .B(CARRYB_19__13_), .CI(SUMB_19__14_), .CO(
        CARRYB_20__13_), .S(SUMB_20__13_) );
  FA_X1 S2_20_14 ( .A(ab_20__14_), .B(CARRYB_19__14_), .CI(SUMB_19__15_), .CO(
        CARRYB_20__14_), .S(SUMB_20__14_) );
  FA_X1 S2_20_15 ( .A(ab_20__15_), .B(CARRYB_19__15_), .CI(SUMB_19__16_), .CO(
        CARRYB_20__15_), .S(SUMB_20__15_) );
  FA_X1 S2_20_16 ( .A(ab_20__16_), .B(CARRYB_19__16_), .CI(SUMB_19__17_), .CO(
        CARRYB_20__16_), .S(SUMB_20__16_) );
  FA_X1 S2_20_17 ( .A(ab_20__17_), .B(CARRYB_19__17_), .CI(SUMB_19__18_), .CO(
        CARRYB_20__17_), .S(SUMB_20__17_) );
  FA_X1 S2_20_18 ( .A(ab_20__18_), .B(CARRYB_19__18_), .CI(SUMB_19__19_), .CO(
        CARRYB_20__18_), .S(SUMB_20__18_) );
  FA_X1 S2_20_19 ( .A(ab_20__19_), .B(CARRYB_19__19_), .CI(SUMB_19__20_), .CO(
        CARRYB_20__19_), .S(SUMB_20__19_) );
  FA_X1 S2_20_20 ( .A(ab_20__20_), .B(CARRYB_19__20_), .CI(SUMB_19__21_), .CO(
        CARRYB_20__20_), .S(SUMB_20__20_) );
  FA_X1 S2_20_21 ( .A(ab_20__21_), .B(CARRYB_19__21_), .CI(SUMB_19__22_), .CO(
        CARRYB_20__21_), .S(SUMB_20__21_) );
  FA_X1 S3_20_22 ( .A(ab_20__22_), .B(CARRYB_19__22_), .CI(A[19]), .CO(
        CARRYB_20__22_), .S(SUMB_20__22_) );
  FA_X1 S1_19_0 ( .A(ab_19__0_), .B(CARRYB_18__0_), .CI(SUMB_18__1_), .CO(
        CARRYB_19__0_), .S(A1_17_) );
  FA_X1 S2_19_1 ( .A(ab_19__1_), .B(CARRYB_18__1_), .CI(SUMB_18__2_), .CO(
        CARRYB_19__1_), .S(SUMB_19__1_) );
  FA_X1 S2_19_2 ( .A(ab_19__2_), .B(CARRYB_18__2_), .CI(SUMB_18__3_), .CO(
        CARRYB_19__2_), .S(SUMB_19__2_) );
  FA_X1 S2_19_3 ( .A(ab_19__3_), .B(CARRYB_18__3_), .CI(SUMB_18__4_), .CO(
        CARRYB_19__3_), .S(SUMB_19__3_) );
  FA_X1 S2_19_4 ( .A(ab_19__4_), .B(CARRYB_18__4_), .CI(SUMB_18__5_), .CO(
        CARRYB_19__4_), .S(SUMB_19__4_) );
  FA_X1 S2_19_5 ( .A(ab_19__5_), .B(CARRYB_18__5_), .CI(SUMB_18__6_), .CO(
        CARRYB_19__5_), .S(SUMB_19__5_) );
  FA_X1 S2_19_6 ( .A(ab_19__6_), .B(CARRYB_18__6_), .CI(SUMB_18__7_), .CO(
        CARRYB_19__6_), .S(SUMB_19__6_) );
  FA_X1 S2_19_7 ( .A(ab_19__7_), .B(CARRYB_18__7_), .CI(SUMB_18__8_), .CO(
        CARRYB_19__7_), .S(SUMB_19__7_) );
  FA_X1 S2_19_8 ( .A(ab_19__8_), .B(CARRYB_18__8_), .CI(SUMB_18__9_), .CO(
        CARRYB_19__8_), .S(SUMB_19__8_) );
  FA_X1 S2_19_9 ( .A(ab_19__9_), .B(CARRYB_18__9_), .CI(SUMB_18__10_), .CO(
        CARRYB_19__9_), .S(SUMB_19__9_) );
  FA_X1 S2_19_10 ( .A(ab_19__10_), .B(CARRYB_18__10_), .CI(SUMB_18__11_), .CO(
        CARRYB_19__10_), .S(SUMB_19__10_) );
  FA_X1 S2_19_11 ( .A(ab_19__11_), .B(CARRYB_18__11_), .CI(SUMB_18__12_), .CO(
        CARRYB_19__11_), .S(SUMB_19__11_) );
  FA_X1 S2_19_12 ( .A(ab_19__12_), .B(CARRYB_18__12_), .CI(SUMB_18__13_), .CO(
        CARRYB_19__12_), .S(SUMB_19__12_) );
  FA_X1 S2_19_13 ( .A(ab_19__13_), .B(CARRYB_18__13_), .CI(SUMB_18__14_), .CO(
        CARRYB_19__13_), .S(SUMB_19__13_) );
  FA_X1 S2_19_14 ( .A(ab_19__14_), .B(CARRYB_18__14_), .CI(SUMB_18__15_), .CO(
        CARRYB_19__14_), .S(SUMB_19__14_) );
  FA_X1 S2_19_15 ( .A(ab_19__15_), .B(CARRYB_18__15_), .CI(SUMB_18__16_), .CO(
        CARRYB_19__15_), .S(SUMB_19__15_) );
  FA_X1 S2_19_16 ( .A(ab_19__16_), .B(CARRYB_18__16_), .CI(SUMB_18__17_), .CO(
        CARRYB_19__16_), .S(SUMB_19__16_) );
  FA_X1 S2_19_17 ( .A(ab_19__17_), .B(CARRYB_18__17_), .CI(SUMB_18__18_), .CO(
        CARRYB_19__17_), .S(SUMB_19__17_) );
  FA_X1 S2_19_18 ( .A(ab_19__18_), .B(CARRYB_18__18_), .CI(SUMB_18__19_), .CO(
        CARRYB_19__18_), .S(SUMB_19__18_) );
  FA_X1 S2_19_19 ( .A(ab_19__19_), .B(CARRYB_18__19_), .CI(SUMB_18__20_), .CO(
        CARRYB_19__19_), .S(SUMB_19__19_) );
  FA_X1 S2_19_20 ( .A(ab_19__20_), .B(CARRYB_18__20_), .CI(SUMB_18__21_), .CO(
        CARRYB_19__20_), .S(SUMB_19__20_) );
  FA_X1 S2_19_21 ( .A(ab_19__21_), .B(CARRYB_18__21_), .CI(SUMB_18__22_), .CO(
        CARRYB_19__21_), .S(SUMB_19__21_) );
  FA_X1 S3_19_22 ( .A(ab_19__22_), .B(CARRYB_18__22_), .CI(A[18]), .CO(
        CARRYB_19__22_), .S(SUMB_19__22_) );
  FA_X1 S1_18_0 ( .A(ab_18__0_), .B(CARRYB_17__0_), .CI(SUMB_17__1_), .CO(
        CARRYB_18__0_), .S(A1_16_) );
  FA_X1 S2_18_1 ( .A(ab_18__1_), .B(CARRYB_17__1_), .CI(SUMB_17__2_), .CO(
        CARRYB_18__1_), .S(SUMB_18__1_) );
  FA_X1 S2_18_2 ( .A(ab_18__2_), .B(CARRYB_17__2_), .CI(SUMB_17__3_), .CO(
        CARRYB_18__2_), .S(SUMB_18__2_) );
  FA_X1 S2_18_3 ( .A(ab_18__3_), .B(CARRYB_17__3_), .CI(SUMB_17__4_), .CO(
        CARRYB_18__3_), .S(SUMB_18__3_) );
  FA_X1 S2_18_4 ( .A(ab_18__4_), .B(CARRYB_17__4_), .CI(SUMB_17__5_), .CO(
        CARRYB_18__4_), .S(SUMB_18__4_) );
  FA_X1 S2_18_5 ( .A(ab_18__5_), .B(CARRYB_17__5_), .CI(SUMB_17__6_), .CO(
        CARRYB_18__5_), .S(SUMB_18__5_) );
  FA_X1 S2_18_6 ( .A(ab_18__6_), .B(CARRYB_17__6_), .CI(SUMB_17__7_), .CO(
        CARRYB_18__6_), .S(SUMB_18__6_) );
  FA_X1 S2_18_7 ( .A(ab_18__7_), .B(CARRYB_17__7_), .CI(SUMB_17__8_), .CO(
        CARRYB_18__7_), .S(SUMB_18__7_) );
  FA_X1 S2_18_8 ( .A(ab_18__8_), .B(CARRYB_17__8_), .CI(SUMB_17__9_), .CO(
        CARRYB_18__8_), .S(SUMB_18__8_) );
  FA_X1 S2_18_9 ( .A(ab_18__9_), .B(CARRYB_17__9_), .CI(SUMB_17__10_), .CO(
        CARRYB_18__9_), .S(SUMB_18__9_) );
  FA_X1 S2_18_10 ( .A(ab_18__10_), .B(CARRYB_17__10_), .CI(SUMB_17__11_), .CO(
        CARRYB_18__10_), .S(SUMB_18__10_) );
  FA_X1 S2_18_11 ( .A(ab_18__11_), .B(CARRYB_17__11_), .CI(SUMB_17__12_), .CO(
        CARRYB_18__11_), .S(SUMB_18__11_) );
  FA_X1 S2_18_12 ( .A(ab_18__12_), .B(CARRYB_17__12_), .CI(SUMB_17__13_), .CO(
        CARRYB_18__12_), .S(SUMB_18__12_) );
  FA_X1 S2_18_13 ( .A(ab_18__13_), .B(CARRYB_17__13_), .CI(SUMB_17__14_), .CO(
        CARRYB_18__13_), .S(SUMB_18__13_) );
  FA_X1 S2_18_14 ( .A(ab_18__14_), .B(CARRYB_17__14_), .CI(SUMB_17__15_), .CO(
        CARRYB_18__14_), .S(SUMB_18__14_) );
  FA_X1 S2_18_15 ( .A(ab_18__15_), .B(CARRYB_17__15_), .CI(SUMB_17__16_), .CO(
        CARRYB_18__15_), .S(SUMB_18__15_) );
  FA_X1 S2_18_16 ( .A(ab_18__16_), .B(CARRYB_17__16_), .CI(SUMB_17__17_), .CO(
        CARRYB_18__16_), .S(SUMB_18__16_) );
  FA_X1 S2_18_17 ( .A(ab_18__17_), .B(CARRYB_17__17_), .CI(SUMB_17__18_), .CO(
        CARRYB_18__17_), .S(SUMB_18__17_) );
  FA_X1 S2_18_18 ( .A(ab_18__18_), .B(CARRYB_17__18_), .CI(SUMB_17__19_), .CO(
        CARRYB_18__18_), .S(SUMB_18__18_) );
  FA_X1 S2_18_19 ( .A(ab_18__19_), .B(CARRYB_17__19_), .CI(SUMB_17__20_), .CO(
        CARRYB_18__19_), .S(SUMB_18__19_) );
  FA_X1 S2_18_20 ( .A(ab_18__20_), .B(CARRYB_17__20_), .CI(SUMB_17__21_), .CO(
        CARRYB_18__20_), .S(SUMB_18__20_) );
  FA_X1 S2_18_21 ( .A(ab_18__21_), .B(CARRYB_17__21_), .CI(SUMB_17__22_), .CO(
        CARRYB_18__21_), .S(SUMB_18__21_) );
  FA_X1 S3_18_22 ( .A(ab_18__22_), .B(CARRYB_17__22_), .CI(A[17]), .CO(
        CARRYB_18__22_), .S(SUMB_18__22_) );
  FA_X1 S1_17_0 ( .A(ab_17__0_), .B(CARRYB_16__0_), .CI(SUMB_16__1_), .CO(
        CARRYB_17__0_), .S(A1_15_) );
  FA_X1 S2_17_1 ( .A(ab_17__1_), .B(CARRYB_16__1_), .CI(SUMB_16__2_), .CO(
        CARRYB_17__1_), .S(SUMB_17__1_) );
  FA_X1 S2_17_2 ( .A(ab_17__2_), .B(CARRYB_16__2_), .CI(SUMB_16__3_), .CO(
        CARRYB_17__2_), .S(SUMB_17__2_) );
  FA_X1 S2_17_3 ( .A(ab_17__3_), .B(CARRYB_16__3_), .CI(SUMB_16__4_), .CO(
        CARRYB_17__3_), .S(SUMB_17__3_) );
  FA_X1 S2_17_4 ( .A(ab_17__4_), .B(CARRYB_16__4_), .CI(SUMB_16__5_), .CO(
        CARRYB_17__4_), .S(SUMB_17__4_) );
  FA_X1 S2_17_5 ( .A(ab_17__5_), .B(CARRYB_16__5_), .CI(SUMB_16__6_), .CO(
        CARRYB_17__5_), .S(SUMB_17__5_) );
  FA_X1 S2_17_6 ( .A(ab_17__6_), .B(CARRYB_16__6_), .CI(SUMB_16__7_), .CO(
        CARRYB_17__6_), .S(SUMB_17__6_) );
  FA_X1 S2_17_7 ( .A(ab_17__7_), .B(CARRYB_16__7_), .CI(SUMB_16__8_), .CO(
        CARRYB_17__7_), .S(SUMB_17__7_) );
  FA_X1 S2_17_8 ( .A(ab_17__8_), .B(CARRYB_16__8_), .CI(SUMB_16__9_), .CO(
        CARRYB_17__8_), .S(SUMB_17__8_) );
  FA_X1 S2_17_9 ( .A(ab_17__9_), .B(CARRYB_16__9_), .CI(SUMB_16__10_), .CO(
        CARRYB_17__9_), .S(SUMB_17__9_) );
  FA_X1 S2_17_10 ( .A(ab_17__10_), .B(CARRYB_16__10_), .CI(SUMB_16__11_), .CO(
        CARRYB_17__10_), .S(SUMB_17__10_) );
  FA_X1 S2_17_11 ( .A(ab_17__11_), .B(CARRYB_16__11_), .CI(SUMB_16__12_), .CO(
        CARRYB_17__11_), .S(SUMB_17__11_) );
  FA_X1 S2_17_12 ( .A(ab_17__12_), .B(CARRYB_16__12_), .CI(SUMB_16__13_), .CO(
        CARRYB_17__12_), .S(SUMB_17__12_) );
  FA_X1 S2_17_13 ( .A(ab_17__13_), .B(CARRYB_16__13_), .CI(SUMB_16__14_), .CO(
        CARRYB_17__13_), .S(SUMB_17__13_) );
  FA_X1 S2_17_14 ( .A(ab_17__14_), .B(CARRYB_16__14_), .CI(SUMB_16__15_), .CO(
        CARRYB_17__14_), .S(SUMB_17__14_) );
  FA_X1 S2_17_15 ( .A(ab_17__15_), .B(CARRYB_16__15_), .CI(SUMB_16__16_), .CO(
        CARRYB_17__15_), .S(SUMB_17__15_) );
  FA_X1 S2_17_16 ( .A(ab_17__16_), .B(CARRYB_16__16_), .CI(SUMB_16__17_), .CO(
        CARRYB_17__16_), .S(SUMB_17__16_) );
  FA_X1 S2_17_17 ( .A(ab_17__17_), .B(CARRYB_16__17_), .CI(SUMB_16__18_), .CO(
        CARRYB_17__17_), .S(SUMB_17__17_) );
  FA_X1 S2_17_18 ( .A(ab_17__18_), .B(CARRYB_16__18_), .CI(SUMB_16__19_), .CO(
        CARRYB_17__18_), .S(SUMB_17__18_) );
  FA_X1 S2_17_19 ( .A(ab_17__19_), .B(CARRYB_16__19_), .CI(SUMB_16__20_), .CO(
        CARRYB_17__19_), .S(SUMB_17__19_) );
  FA_X1 S2_17_20 ( .A(ab_17__20_), .B(CARRYB_16__20_), .CI(SUMB_16__21_), .CO(
        CARRYB_17__20_), .S(SUMB_17__20_) );
  FA_X1 S2_17_21 ( .A(ab_17__21_), .B(CARRYB_16__21_), .CI(SUMB_16__22_), .CO(
        CARRYB_17__21_), .S(SUMB_17__21_) );
  FA_X1 S3_17_22 ( .A(ab_17__22_), .B(CARRYB_16__22_), .CI(A[16]), .CO(
        CARRYB_17__22_), .S(SUMB_17__22_) );
  FA_X1 S1_16_0 ( .A(ab_16__0_), .B(CARRYB_15__0_), .CI(SUMB_15__1_), .CO(
        CARRYB_16__0_), .S(A1_14_) );
  FA_X1 S2_16_1 ( .A(ab_16__1_), .B(CARRYB_15__1_), .CI(SUMB_15__2_), .CO(
        CARRYB_16__1_), .S(SUMB_16__1_) );
  FA_X1 S2_16_2 ( .A(ab_16__2_), .B(CARRYB_15__2_), .CI(SUMB_15__3_), .CO(
        CARRYB_16__2_), .S(SUMB_16__2_) );
  FA_X1 S2_16_3 ( .A(ab_16__3_), .B(CARRYB_15__3_), .CI(SUMB_15__4_), .CO(
        CARRYB_16__3_), .S(SUMB_16__3_) );
  FA_X1 S2_16_4 ( .A(ab_16__4_), .B(CARRYB_15__4_), .CI(SUMB_15__5_), .CO(
        CARRYB_16__4_), .S(SUMB_16__4_) );
  FA_X1 S2_16_5 ( .A(ab_16__5_), .B(CARRYB_15__5_), .CI(SUMB_15__6_), .CO(
        CARRYB_16__5_), .S(SUMB_16__5_) );
  FA_X1 S2_16_6 ( .A(ab_16__6_), .B(CARRYB_15__6_), .CI(SUMB_15__7_), .CO(
        CARRYB_16__6_), .S(SUMB_16__6_) );
  FA_X1 S2_16_7 ( .A(ab_16__7_), .B(CARRYB_15__7_), .CI(SUMB_15__8_), .CO(
        CARRYB_16__7_), .S(SUMB_16__7_) );
  FA_X1 S2_16_8 ( .A(ab_16__8_), .B(CARRYB_15__8_), .CI(SUMB_15__9_), .CO(
        CARRYB_16__8_), .S(SUMB_16__8_) );
  FA_X1 S2_16_9 ( .A(ab_16__9_), .B(CARRYB_15__9_), .CI(SUMB_15__10_), .CO(
        CARRYB_16__9_), .S(SUMB_16__9_) );
  FA_X1 S2_16_10 ( .A(ab_16__10_), .B(CARRYB_15__10_), .CI(SUMB_15__11_), .CO(
        CARRYB_16__10_), .S(SUMB_16__10_) );
  FA_X1 S2_16_11 ( .A(ab_16__11_), .B(CARRYB_15__11_), .CI(SUMB_15__12_), .CO(
        CARRYB_16__11_), .S(SUMB_16__11_) );
  FA_X1 S2_16_12 ( .A(ab_16__12_), .B(CARRYB_15__12_), .CI(SUMB_15__13_), .CO(
        CARRYB_16__12_), .S(SUMB_16__12_) );
  FA_X1 S2_16_13 ( .A(ab_16__13_), .B(CARRYB_15__13_), .CI(SUMB_15__14_), .CO(
        CARRYB_16__13_), .S(SUMB_16__13_) );
  FA_X1 S2_16_14 ( .A(ab_16__14_), .B(CARRYB_15__14_), .CI(SUMB_15__15_), .CO(
        CARRYB_16__14_), .S(SUMB_16__14_) );
  FA_X1 S2_16_15 ( .A(ab_16__15_), .B(CARRYB_15__15_), .CI(SUMB_15__16_), .CO(
        CARRYB_16__15_), .S(SUMB_16__15_) );
  FA_X1 S2_16_16 ( .A(ab_16__16_), .B(CARRYB_15__16_), .CI(SUMB_15__17_), .CO(
        CARRYB_16__16_), .S(SUMB_16__16_) );
  FA_X1 S2_16_17 ( .A(ab_16__17_), .B(CARRYB_15__17_), .CI(SUMB_15__18_), .CO(
        CARRYB_16__17_), .S(SUMB_16__17_) );
  FA_X1 S2_16_18 ( .A(ab_16__18_), .B(CARRYB_15__18_), .CI(SUMB_15__19_), .CO(
        CARRYB_16__18_), .S(SUMB_16__18_) );
  FA_X1 S2_16_19 ( .A(ab_16__19_), .B(CARRYB_15__19_), .CI(SUMB_15__20_), .CO(
        CARRYB_16__19_), .S(SUMB_16__19_) );
  FA_X1 S2_16_20 ( .A(ab_16__20_), .B(CARRYB_15__20_), .CI(SUMB_15__21_), .CO(
        CARRYB_16__20_), .S(SUMB_16__20_) );
  FA_X1 S2_16_21 ( .A(ab_16__21_), .B(CARRYB_15__21_), .CI(SUMB_15__22_), .CO(
        CARRYB_16__21_), .S(SUMB_16__21_) );
  FA_X1 S3_16_22 ( .A(ab_16__22_), .B(CARRYB_15__22_), .CI(A[15]), .CO(
        CARRYB_16__22_), .S(SUMB_16__22_) );
  FA_X1 S1_15_0 ( .A(ab_15__0_), .B(CARRYB_14__0_), .CI(SUMB_14__1_), .CO(
        CARRYB_15__0_), .S(A1_13_) );
  FA_X1 S2_15_1 ( .A(ab_15__1_), .B(CARRYB_14__1_), .CI(SUMB_14__2_), .CO(
        CARRYB_15__1_), .S(SUMB_15__1_) );
  FA_X1 S2_15_2 ( .A(ab_15__2_), .B(CARRYB_14__2_), .CI(SUMB_14__3_), .CO(
        CARRYB_15__2_), .S(SUMB_15__2_) );
  FA_X1 S2_15_3 ( .A(ab_15__3_), .B(CARRYB_14__3_), .CI(SUMB_14__4_), .CO(
        CARRYB_15__3_), .S(SUMB_15__3_) );
  FA_X1 S2_15_4 ( .A(ab_15__4_), .B(CARRYB_14__4_), .CI(SUMB_14__5_), .CO(
        CARRYB_15__4_), .S(SUMB_15__4_) );
  FA_X1 S2_15_5 ( .A(ab_15__5_), .B(CARRYB_14__5_), .CI(SUMB_14__6_), .CO(
        CARRYB_15__5_), .S(SUMB_15__5_) );
  FA_X1 S2_15_6 ( .A(ab_15__6_), .B(CARRYB_14__6_), .CI(SUMB_14__7_), .CO(
        CARRYB_15__6_), .S(SUMB_15__6_) );
  FA_X1 S2_15_7 ( .A(ab_15__7_), .B(CARRYB_14__7_), .CI(SUMB_14__8_), .CO(
        CARRYB_15__7_), .S(SUMB_15__7_) );
  FA_X1 S2_15_8 ( .A(ab_15__8_), .B(CARRYB_14__8_), .CI(SUMB_14__9_), .CO(
        CARRYB_15__8_), .S(SUMB_15__8_) );
  FA_X1 S2_15_9 ( .A(ab_15__9_), .B(CARRYB_14__9_), .CI(SUMB_14__10_), .CO(
        CARRYB_15__9_), .S(SUMB_15__9_) );
  FA_X1 S2_15_10 ( .A(ab_15__10_), .B(CARRYB_14__10_), .CI(SUMB_14__11_), .CO(
        CARRYB_15__10_), .S(SUMB_15__10_) );
  FA_X1 S2_15_11 ( .A(ab_15__11_), .B(CARRYB_14__11_), .CI(SUMB_14__12_), .CO(
        CARRYB_15__11_), .S(SUMB_15__11_) );
  FA_X1 S2_15_12 ( .A(ab_15__12_), .B(CARRYB_14__12_), .CI(SUMB_14__13_), .CO(
        CARRYB_15__12_), .S(SUMB_15__12_) );
  FA_X1 S2_15_13 ( .A(ab_15__13_), .B(CARRYB_14__13_), .CI(SUMB_14__14_), .CO(
        CARRYB_15__13_), .S(SUMB_15__13_) );
  FA_X1 S2_15_14 ( .A(ab_15__14_), .B(CARRYB_14__14_), .CI(SUMB_14__15_), .CO(
        CARRYB_15__14_), .S(SUMB_15__14_) );
  FA_X1 S2_15_15 ( .A(ab_15__15_), .B(CARRYB_14__15_), .CI(SUMB_14__16_), .CO(
        CARRYB_15__15_), .S(SUMB_15__15_) );
  FA_X1 S2_15_16 ( .A(ab_15__16_), .B(CARRYB_14__16_), .CI(SUMB_14__17_), .CO(
        CARRYB_15__16_), .S(SUMB_15__16_) );
  FA_X1 S2_15_17 ( .A(ab_15__17_), .B(CARRYB_14__17_), .CI(SUMB_14__18_), .CO(
        CARRYB_15__17_), .S(SUMB_15__17_) );
  FA_X1 S2_15_18 ( .A(ab_15__18_), .B(CARRYB_14__18_), .CI(SUMB_14__19_), .CO(
        CARRYB_15__18_), .S(SUMB_15__18_) );
  FA_X1 S2_15_19 ( .A(ab_15__19_), .B(CARRYB_14__19_), .CI(SUMB_14__20_), .CO(
        CARRYB_15__19_), .S(SUMB_15__19_) );
  FA_X1 S2_15_20 ( .A(ab_15__20_), .B(CARRYB_14__20_), .CI(SUMB_14__21_), .CO(
        CARRYB_15__20_), .S(SUMB_15__20_) );
  FA_X1 S2_15_21 ( .A(ab_15__21_), .B(CARRYB_14__21_), .CI(SUMB_14__22_), .CO(
        CARRYB_15__21_), .S(SUMB_15__21_) );
  FA_X1 S3_15_22 ( .A(ab_15__22_), .B(CARRYB_14__22_), .CI(A[14]), .CO(
        CARRYB_15__22_), .S(SUMB_15__22_) );
  FA_X1 S1_14_0 ( .A(ab_14__0_), .B(CARRYB_13__0_), .CI(SUMB_13__1_), .CO(
        CARRYB_14__0_), .S(A1_12_) );
  FA_X1 S2_14_1 ( .A(ab_14__1_), .B(CARRYB_13__1_), .CI(SUMB_13__2_), .CO(
        CARRYB_14__1_), .S(SUMB_14__1_) );
  FA_X1 S2_14_2 ( .A(ab_14__2_), .B(CARRYB_13__2_), .CI(SUMB_13__3_), .CO(
        CARRYB_14__2_), .S(SUMB_14__2_) );
  FA_X1 S2_14_3 ( .A(ab_14__3_), .B(CARRYB_13__3_), .CI(SUMB_13__4_), .CO(
        CARRYB_14__3_), .S(SUMB_14__3_) );
  FA_X1 S2_14_4 ( .A(ab_14__4_), .B(CARRYB_13__4_), .CI(SUMB_13__5_), .CO(
        CARRYB_14__4_), .S(SUMB_14__4_) );
  FA_X1 S2_14_5 ( .A(ab_14__5_), .B(CARRYB_13__5_), .CI(SUMB_13__6_), .CO(
        CARRYB_14__5_), .S(SUMB_14__5_) );
  FA_X1 S2_14_6 ( .A(ab_14__6_), .B(CARRYB_13__6_), .CI(SUMB_13__7_), .CO(
        CARRYB_14__6_), .S(SUMB_14__6_) );
  FA_X1 S2_14_7 ( .A(ab_14__7_), .B(CARRYB_13__7_), .CI(SUMB_13__8_), .CO(
        CARRYB_14__7_), .S(SUMB_14__7_) );
  FA_X1 S2_14_8 ( .A(ab_14__8_), .B(CARRYB_13__8_), .CI(SUMB_13__9_), .CO(
        CARRYB_14__8_), .S(SUMB_14__8_) );
  FA_X1 S2_14_9 ( .A(ab_14__9_), .B(CARRYB_13__9_), .CI(SUMB_13__10_), .CO(
        CARRYB_14__9_), .S(SUMB_14__9_) );
  FA_X1 S2_14_10 ( .A(ab_14__10_), .B(CARRYB_13__10_), .CI(SUMB_13__11_), .CO(
        CARRYB_14__10_), .S(SUMB_14__10_) );
  FA_X1 S2_14_11 ( .A(ab_14__11_), .B(CARRYB_13__11_), .CI(SUMB_13__12_), .CO(
        CARRYB_14__11_), .S(SUMB_14__11_) );
  FA_X1 S2_14_12 ( .A(ab_14__12_), .B(CARRYB_13__12_), .CI(SUMB_13__13_), .CO(
        CARRYB_14__12_), .S(SUMB_14__12_) );
  FA_X1 S2_14_13 ( .A(ab_14__13_), .B(CARRYB_13__13_), .CI(SUMB_13__14_), .CO(
        CARRYB_14__13_), .S(SUMB_14__13_) );
  FA_X1 S2_14_14 ( .A(ab_14__14_), .B(CARRYB_13__14_), .CI(SUMB_13__15_), .CO(
        CARRYB_14__14_), .S(SUMB_14__14_) );
  FA_X1 S2_14_15 ( .A(ab_14__15_), .B(CARRYB_13__15_), .CI(SUMB_13__16_), .CO(
        CARRYB_14__15_), .S(SUMB_14__15_) );
  FA_X1 S2_14_16 ( .A(ab_14__16_), .B(CARRYB_13__16_), .CI(SUMB_13__17_), .CO(
        CARRYB_14__16_), .S(SUMB_14__16_) );
  FA_X1 S2_14_17 ( .A(ab_14__17_), .B(CARRYB_13__17_), .CI(SUMB_13__18_), .CO(
        CARRYB_14__17_), .S(SUMB_14__17_) );
  FA_X1 S2_14_18 ( .A(ab_14__18_), .B(CARRYB_13__18_), .CI(SUMB_13__19_), .CO(
        CARRYB_14__18_), .S(SUMB_14__18_) );
  FA_X1 S2_14_19 ( .A(ab_14__19_), .B(CARRYB_13__19_), .CI(SUMB_13__20_), .CO(
        CARRYB_14__19_), .S(SUMB_14__19_) );
  FA_X1 S2_14_20 ( .A(ab_14__20_), .B(CARRYB_13__20_), .CI(SUMB_13__21_), .CO(
        CARRYB_14__20_), .S(SUMB_14__20_) );
  FA_X1 S2_14_21 ( .A(ab_14__21_), .B(CARRYB_13__21_), .CI(SUMB_13__22_), .CO(
        CARRYB_14__21_), .S(SUMB_14__21_) );
  FA_X1 S3_14_22 ( .A(ab_14__22_), .B(CARRYB_13__22_), .CI(A[13]), .CO(
        CARRYB_14__22_), .S(SUMB_14__22_) );
  FA_X1 S1_13_0 ( .A(ab_13__0_), .B(CARRYB_12__0_), .CI(SUMB_12__1_), .CO(
        CARRYB_13__0_), .S(A1_11_) );
  FA_X1 S2_13_1 ( .A(ab_13__1_), .B(CARRYB_12__1_), .CI(SUMB_12__2_), .CO(
        CARRYB_13__1_), .S(SUMB_13__1_) );
  FA_X1 S2_13_2 ( .A(ab_13__2_), .B(CARRYB_12__2_), .CI(SUMB_12__3_), .CO(
        CARRYB_13__2_), .S(SUMB_13__2_) );
  FA_X1 S2_13_3 ( .A(ab_13__3_), .B(CARRYB_12__3_), .CI(SUMB_12__4_), .CO(
        CARRYB_13__3_), .S(SUMB_13__3_) );
  FA_X1 S2_13_4 ( .A(ab_13__4_), .B(CARRYB_12__4_), .CI(SUMB_12__5_), .CO(
        CARRYB_13__4_), .S(SUMB_13__4_) );
  FA_X1 S2_13_5 ( .A(ab_13__5_), .B(CARRYB_12__5_), .CI(SUMB_12__6_), .CO(
        CARRYB_13__5_), .S(SUMB_13__5_) );
  FA_X1 S2_13_6 ( .A(ab_13__6_), .B(CARRYB_12__6_), .CI(SUMB_12__7_), .CO(
        CARRYB_13__6_), .S(SUMB_13__6_) );
  FA_X1 S2_13_7 ( .A(ab_13__7_), .B(CARRYB_12__7_), .CI(SUMB_12__8_), .CO(
        CARRYB_13__7_), .S(SUMB_13__7_) );
  FA_X1 S2_13_8 ( .A(ab_13__8_), .B(CARRYB_12__8_), .CI(SUMB_12__9_), .CO(
        CARRYB_13__8_), .S(SUMB_13__8_) );
  FA_X1 S2_13_9 ( .A(ab_13__9_), .B(CARRYB_12__9_), .CI(SUMB_12__10_), .CO(
        CARRYB_13__9_), .S(SUMB_13__9_) );
  FA_X1 S2_13_10 ( .A(ab_13__10_), .B(CARRYB_12__10_), .CI(SUMB_12__11_), .CO(
        CARRYB_13__10_), .S(SUMB_13__10_) );
  FA_X1 S2_13_11 ( .A(ab_13__11_), .B(CARRYB_12__11_), .CI(SUMB_12__12_), .CO(
        CARRYB_13__11_), .S(SUMB_13__11_) );
  FA_X1 S2_13_12 ( .A(ab_13__12_), .B(CARRYB_12__12_), .CI(SUMB_12__13_), .CO(
        CARRYB_13__12_), .S(SUMB_13__12_) );
  FA_X1 S2_13_13 ( .A(ab_13__13_), .B(CARRYB_12__13_), .CI(SUMB_12__14_), .CO(
        CARRYB_13__13_), .S(SUMB_13__13_) );
  FA_X1 S2_13_14 ( .A(ab_13__14_), .B(CARRYB_12__14_), .CI(SUMB_12__15_), .CO(
        CARRYB_13__14_), .S(SUMB_13__14_) );
  FA_X1 S2_13_15 ( .A(ab_13__15_), .B(CARRYB_12__15_), .CI(SUMB_12__16_), .CO(
        CARRYB_13__15_), .S(SUMB_13__15_) );
  FA_X1 S2_13_16 ( .A(ab_13__16_), .B(CARRYB_12__16_), .CI(SUMB_12__17_), .CO(
        CARRYB_13__16_), .S(SUMB_13__16_) );
  FA_X1 S2_13_17 ( .A(ab_13__17_), .B(CARRYB_12__17_), .CI(SUMB_12__18_), .CO(
        CARRYB_13__17_), .S(SUMB_13__17_) );
  FA_X1 S2_13_18 ( .A(ab_13__18_), .B(CARRYB_12__18_), .CI(SUMB_12__19_), .CO(
        CARRYB_13__18_), .S(SUMB_13__18_) );
  FA_X1 S2_13_19 ( .A(ab_13__19_), .B(CARRYB_12__19_), .CI(SUMB_12__20_), .CO(
        CARRYB_13__19_), .S(SUMB_13__19_) );
  FA_X1 S2_13_20 ( .A(ab_13__20_), .B(CARRYB_12__20_), .CI(SUMB_12__21_), .CO(
        CARRYB_13__20_), .S(SUMB_13__20_) );
  FA_X1 S2_13_21 ( .A(ab_13__21_), .B(CARRYB_12__21_), .CI(SUMB_12__22_), .CO(
        CARRYB_13__21_), .S(SUMB_13__21_) );
  FA_X1 S3_13_22 ( .A(ab_13__22_), .B(CARRYB_12__22_), .CI(A[12]), .CO(
        CARRYB_13__22_), .S(SUMB_13__22_) );
  FA_X1 S1_12_0 ( .A(ab_12__0_), .B(CARRYB_11__0_), .CI(SUMB_11__1_), .CO(
        CARRYB_12__0_), .S(A1_10_) );
  FA_X1 S2_12_1 ( .A(ab_12__1_), .B(CARRYB_11__1_), .CI(SUMB_11__2_), .CO(
        CARRYB_12__1_), .S(SUMB_12__1_) );
  FA_X1 S2_12_2 ( .A(ab_12__2_), .B(CARRYB_11__2_), .CI(SUMB_11__3_), .CO(
        CARRYB_12__2_), .S(SUMB_12__2_) );
  FA_X1 S2_12_3 ( .A(ab_12__3_), .B(CARRYB_11__3_), .CI(SUMB_11__4_), .CO(
        CARRYB_12__3_), .S(SUMB_12__3_) );
  FA_X1 S2_12_4 ( .A(ab_12__4_), .B(CARRYB_11__4_), .CI(SUMB_11__5_), .CO(
        CARRYB_12__4_), .S(SUMB_12__4_) );
  FA_X1 S2_12_5 ( .A(ab_12__5_), .B(CARRYB_11__5_), .CI(SUMB_11__6_), .CO(
        CARRYB_12__5_), .S(SUMB_12__5_) );
  FA_X1 S2_12_6 ( .A(ab_12__6_), .B(CARRYB_11__6_), .CI(SUMB_11__7_), .CO(
        CARRYB_12__6_), .S(SUMB_12__6_) );
  FA_X1 S2_12_7 ( .A(ab_12__7_), .B(CARRYB_11__7_), .CI(SUMB_11__8_), .CO(
        CARRYB_12__7_), .S(SUMB_12__7_) );
  FA_X1 S2_12_8 ( .A(ab_12__8_), .B(CARRYB_11__8_), .CI(SUMB_11__9_), .CO(
        CARRYB_12__8_), .S(SUMB_12__8_) );
  FA_X1 S2_12_9 ( .A(ab_12__9_), .B(CARRYB_11__9_), .CI(SUMB_11__10_), .CO(
        CARRYB_12__9_), .S(SUMB_12__9_) );
  FA_X1 S2_12_10 ( .A(ab_12__10_), .B(CARRYB_11__10_), .CI(SUMB_11__11_), .CO(
        CARRYB_12__10_), .S(SUMB_12__10_) );
  FA_X1 S2_12_11 ( .A(ab_12__11_), .B(CARRYB_11__11_), .CI(SUMB_11__12_), .CO(
        CARRYB_12__11_), .S(SUMB_12__11_) );
  FA_X1 S2_12_12 ( .A(ab_12__12_), .B(CARRYB_11__12_), .CI(SUMB_11__13_), .CO(
        CARRYB_12__12_), .S(SUMB_12__12_) );
  FA_X1 S2_12_13 ( .A(ab_12__13_), .B(CARRYB_11__13_), .CI(SUMB_11__14_), .CO(
        CARRYB_12__13_), .S(SUMB_12__13_) );
  FA_X1 S2_12_14 ( .A(ab_12__14_), .B(CARRYB_11__14_), .CI(SUMB_11__15_), .CO(
        CARRYB_12__14_), .S(SUMB_12__14_) );
  FA_X1 S2_12_15 ( .A(ab_12__15_), .B(CARRYB_11__15_), .CI(SUMB_11__16_), .CO(
        CARRYB_12__15_), .S(SUMB_12__15_) );
  FA_X1 S2_12_16 ( .A(ab_12__16_), .B(CARRYB_11__16_), .CI(SUMB_11__17_), .CO(
        CARRYB_12__16_), .S(SUMB_12__16_) );
  FA_X1 S2_12_17 ( .A(ab_12__17_), .B(CARRYB_11__17_), .CI(SUMB_11__18_), .CO(
        CARRYB_12__17_), .S(SUMB_12__17_) );
  FA_X1 S2_12_18 ( .A(ab_12__18_), .B(CARRYB_11__18_), .CI(SUMB_11__19_), .CO(
        CARRYB_12__18_), .S(SUMB_12__18_) );
  FA_X1 S2_12_19 ( .A(ab_12__19_), .B(CARRYB_11__19_), .CI(SUMB_11__20_), .CO(
        CARRYB_12__19_), .S(SUMB_12__19_) );
  FA_X1 S2_12_20 ( .A(ab_12__20_), .B(CARRYB_11__20_), .CI(SUMB_11__21_), .CO(
        CARRYB_12__20_), .S(SUMB_12__20_) );
  FA_X1 S2_12_21 ( .A(ab_12__21_), .B(CARRYB_11__21_), .CI(SUMB_11__22_), .CO(
        CARRYB_12__21_), .S(SUMB_12__21_) );
  FA_X1 S3_12_22 ( .A(ab_12__22_), .B(CARRYB_11__22_), .CI(A[11]), .CO(
        CARRYB_12__22_), .S(SUMB_12__22_) );
  FA_X1 S1_11_0 ( .A(ab_11__0_), .B(CARRYB_10__0_), .CI(SUMB_10__1_), .CO(
        CARRYB_11__0_), .S(A1_9_) );
  FA_X1 S2_11_1 ( .A(ab_11__1_), .B(CARRYB_10__1_), .CI(SUMB_10__2_), .CO(
        CARRYB_11__1_), .S(SUMB_11__1_) );
  FA_X1 S2_11_2 ( .A(ab_11__2_), .B(CARRYB_10__2_), .CI(SUMB_10__3_), .CO(
        CARRYB_11__2_), .S(SUMB_11__2_) );
  FA_X1 S2_11_3 ( .A(ab_11__3_), .B(CARRYB_10__3_), .CI(SUMB_10__4_), .CO(
        CARRYB_11__3_), .S(SUMB_11__3_) );
  FA_X1 S2_11_4 ( .A(ab_11__4_), .B(CARRYB_10__4_), .CI(SUMB_10__5_), .CO(
        CARRYB_11__4_), .S(SUMB_11__4_) );
  FA_X1 S2_11_5 ( .A(ab_11__5_), .B(CARRYB_10__5_), .CI(SUMB_10__6_), .CO(
        CARRYB_11__5_), .S(SUMB_11__5_) );
  FA_X1 S2_11_6 ( .A(ab_11__6_), .B(CARRYB_10__6_), .CI(SUMB_10__7_), .CO(
        CARRYB_11__6_), .S(SUMB_11__6_) );
  FA_X1 S2_11_7 ( .A(ab_11__7_), .B(CARRYB_10__7_), .CI(SUMB_10__8_), .CO(
        CARRYB_11__7_), .S(SUMB_11__7_) );
  FA_X1 S2_11_8 ( .A(ab_11__8_), .B(CARRYB_10__8_), .CI(SUMB_10__9_), .CO(
        CARRYB_11__8_), .S(SUMB_11__8_) );
  FA_X1 S2_11_9 ( .A(ab_11__9_), .B(CARRYB_10__9_), .CI(SUMB_10__10_), .CO(
        CARRYB_11__9_), .S(SUMB_11__9_) );
  FA_X1 S2_11_10 ( .A(ab_11__10_), .B(CARRYB_10__10_), .CI(SUMB_10__11_), .CO(
        CARRYB_11__10_), .S(SUMB_11__10_) );
  FA_X1 S2_11_11 ( .A(ab_11__11_), .B(CARRYB_10__11_), .CI(SUMB_10__12_), .CO(
        CARRYB_11__11_), .S(SUMB_11__11_) );
  FA_X1 S2_11_12 ( .A(ab_11__12_), .B(CARRYB_10__12_), .CI(SUMB_10__13_), .CO(
        CARRYB_11__12_), .S(SUMB_11__12_) );
  FA_X1 S2_11_13 ( .A(ab_11__13_), .B(CARRYB_10__13_), .CI(SUMB_10__14_), .CO(
        CARRYB_11__13_), .S(SUMB_11__13_) );
  FA_X1 S2_11_14 ( .A(ab_11__14_), .B(CARRYB_10__14_), .CI(SUMB_10__15_), .CO(
        CARRYB_11__14_), .S(SUMB_11__14_) );
  FA_X1 S2_11_15 ( .A(ab_11__15_), .B(CARRYB_10__15_), .CI(SUMB_10__16_), .CO(
        CARRYB_11__15_), .S(SUMB_11__15_) );
  FA_X1 S2_11_16 ( .A(ab_11__16_), .B(CARRYB_10__16_), .CI(SUMB_10__17_), .CO(
        CARRYB_11__16_), .S(SUMB_11__16_) );
  FA_X1 S2_11_17 ( .A(ab_11__17_), .B(CARRYB_10__17_), .CI(SUMB_10__18_), .CO(
        CARRYB_11__17_), .S(SUMB_11__17_) );
  FA_X1 S2_11_18 ( .A(ab_11__18_), .B(CARRYB_10__18_), .CI(SUMB_10__19_), .CO(
        CARRYB_11__18_), .S(SUMB_11__18_) );
  FA_X1 S2_11_19 ( .A(ab_11__19_), .B(CARRYB_10__19_), .CI(SUMB_10__20_), .CO(
        CARRYB_11__19_), .S(SUMB_11__19_) );
  FA_X1 S2_11_20 ( .A(ab_11__20_), .B(CARRYB_10__20_), .CI(SUMB_10__21_), .CO(
        CARRYB_11__20_), .S(SUMB_11__20_) );
  FA_X1 S2_11_21 ( .A(ab_11__21_), .B(CARRYB_10__21_), .CI(SUMB_10__22_), .CO(
        CARRYB_11__21_), .S(SUMB_11__21_) );
  FA_X1 S3_11_22 ( .A(ab_11__22_), .B(CARRYB_10__22_), .CI(A[10]), .CO(
        CARRYB_11__22_), .S(SUMB_11__22_) );
  FA_X1 S1_10_0 ( .A(ab_10__0_), .B(CARRYB_9__0_), .CI(SUMB_9__1_), .CO(
        CARRYB_10__0_), .S(A1_8_) );
  FA_X1 S2_10_1 ( .A(ab_10__1_), .B(CARRYB_9__1_), .CI(SUMB_9__2_), .CO(
        CARRYB_10__1_), .S(SUMB_10__1_) );
  FA_X1 S2_10_2 ( .A(ab_10__2_), .B(CARRYB_9__2_), .CI(SUMB_9__3_), .CO(
        CARRYB_10__2_), .S(SUMB_10__2_) );
  FA_X1 S2_10_3 ( .A(ab_10__3_), .B(CARRYB_9__3_), .CI(SUMB_9__4_), .CO(
        CARRYB_10__3_), .S(SUMB_10__3_) );
  FA_X1 S2_10_4 ( .A(ab_10__4_), .B(CARRYB_9__4_), .CI(SUMB_9__5_), .CO(
        CARRYB_10__4_), .S(SUMB_10__4_) );
  FA_X1 S2_10_5 ( .A(ab_10__5_), .B(CARRYB_9__5_), .CI(SUMB_9__6_), .CO(
        CARRYB_10__5_), .S(SUMB_10__5_) );
  FA_X1 S2_10_6 ( .A(ab_10__6_), .B(CARRYB_9__6_), .CI(SUMB_9__7_), .CO(
        CARRYB_10__6_), .S(SUMB_10__6_) );
  FA_X1 S2_10_7 ( .A(ab_10__7_), .B(CARRYB_9__7_), .CI(SUMB_9__8_), .CO(
        CARRYB_10__7_), .S(SUMB_10__7_) );
  FA_X1 S2_10_8 ( .A(ab_10__8_), .B(CARRYB_9__8_), .CI(SUMB_9__9_), .CO(
        CARRYB_10__8_), .S(SUMB_10__8_) );
  FA_X1 S2_10_9 ( .A(ab_10__9_), .B(CARRYB_9__9_), .CI(SUMB_9__10_), .CO(
        CARRYB_10__9_), .S(SUMB_10__9_) );
  FA_X1 S2_10_10 ( .A(ab_10__10_), .B(CARRYB_9__10_), .CI(SUMB_9__11_), .CO(
        CARRYB_10__10_), .S(SUMB_10__10_) );
  FA_X1 S2_10_11 ( .A(ab_10__11_), .B(CARRYB_9__11_), .CI(SUMB_9__12_), .CO(
        CARRYB_10__11_), .S(SUMB_10__11_) );
  FA_X1 S2_10_12 ( .A(ab_10__12_), .B(CARRYB_9__12_), .CI(SUMB_9__13_), .CO(
        CARRYB_10__12_), .S(SUMB_10__12_) );
  FA_X1 S2_10_13 ( .A(ab_10__13_), .B(CARRYB_9__13_), .CI(SUMB_9__14_), .CO(
        CARRYB_10__13_), .S(SUMB_10__13_) );
  FA_X1 S2_10_14 ( .A(ab_10__14_), .B(CARRYB_9__14_), .CI(SUMB_9__15_), .CO(
        CARRYB_10__14_), .S(SUMB_10__14_) );
  FA_X1 S2_10_15 ( .A(ab_10__15_), .B(CARRYB_9__15_), .CI(SUMB_9__16_), .CO(
        CARRYB_10__15_), .S(SUMB_10__15_) );
  FA_X1 S2_10_16 ( .A(ab_10__16_), .B(CARRYB_9__16_), .CI(SUMB_9__17_), .CO(
        CARRYB_10__16_), .S(SUMB_10__16_) );
  FA_X1 S2_10_17 ( .A(ab_10__17_), .B(CARRYB_9__17_), .CI(SUMB_9__18_), .CO(
        CARRYB_10__17_), .S(SUMB_10__17_) );
  FA_X1 S2_10_18 ( .A(ab_10__18_), .B(CARRYB_9__18_), .CI(SUMB_9__19_), .CO(
        CARRYB_10__18_), .S(SUMB_10__18_) );
  FA_X1 S2_10_19 ( .A(ab_10__19_), .B(CARRYB_9__19_), .CI(SUMB_9__20_), .CO(
        CARRYB_10__19_), .S(SUMB_10__19_) );
  FA_X1 S2_10_20 ( .A(ab_10__20_), .B(CARRYB_9__20_), .CI(SUMB_9__21_), .CO(
        CARRYB_10__20_), .S(SUMB_10__20_) );
  FA_X1 S2_10_21 ( .A(ab_10__21_), .B(CARRYB_9__21_), .CI(SUMB_9__22_), .CO(
        CARRYB_10__21_), .S(SUMB_10__21_) );
  FA_X1 S3_10_22 ( .A(ab_10__22_), .B(CARRYB_9__22_), .CI(A[9]), .CO(
        CARRYB_10__22_), .S(SUMB_10__22_) );
  FA_X1 S1_9_0 ( .A(ab_9__0_), .B(CARRYB_8__0_), .CI(SUMB_8__1_), .CO(
        CARRYB_9__0_), .S(A1_7_) );
  FA_X1 S2_9_1 ( .A(ab_9__1_), .B(CARRYB_8__1_), .CI(SUMB_8__2_), .CO(
        CARRYB_9__1_), .S(SUMB_9__1_) );
  FA_X1 S2_9_2 ( .A(ab_9__2_), .B(CARRYB_8__2_), .CI(SUMB_8__3_), .CO(
        CARRYB_9__2_), .S(SUMB_9__2_) );
  FA_X1 S2_9_3 ( .A(ab_9__3_), .B(CARRYB_8__3_), .CI(SUMB_8__4_), .CO(
        CARRYB_9__3_), .S(SUMB_9__3_) );
  FA_X1 S2_9_4 ( .A(ab_9__4_), .B(CARRYB_8__4_), .CI(SUMB_8__5_), .CO(
        CARRYB_9__4_), .S(SUMB_9__4_) );
  FA_X1 S2_9_5 ( .A(ab_9__5_), .B(CARRYB_8__5_), .CI(SUMB_8__6_), .CO(
        CARRYB_9__5_), .S(SUMB_9__5_) );
  FA_X1 S2_9_6 ( .A(ab_9__6_), .B(CARRYB_8__6_), .CI(SUMB_8__7_), .CO(
        CARRYB_9__6_), .S(SUMB_9__6_) );
  FA_X1 S2_9_7 ( .A(ab_9__7_), .B(CARRYB_8__7_), .CI(SUMB_8__8_), .CO(
        CARRYB_9__7_), .S(SUMB_9__7_) );
  FA_X1 S2_9_8 ( .A(ab_9__8_), .B(CARRYB_8__8_), .CI(SUMB_8__9_), .CO(
        CARRYB_9__8_), .S(SUMB_9__8_) );
  FA_X1 S2_9_9 ( .A(ab_9__9_), .B(CARRYB_8__9_), .CI(SUMB_8__10_), .CO(
        CARRYB_9__9_), .S(SUMB_9__9_) );
  FA_X1 S2_9_10 ( .A(ab_9__10_), .B(CARRYB_8__10_), .CI(SUMB_8__11_), .CO(
        CARRYB_9__10_), .S(SUMB_9__10_) );
  FA_X1 S2_9_11 ( .A(ab_9__11_), .B(CARRYB_8__11_), .CI(SUMB_8__12_), .CO(
        CARRYB_9__11_), .S(SUMB_9__11_) );
  FA_X1 S2_9_12 ( .A(ab_9__12_), .B(CARRYB_8__12_), .CI(SUMB_8__13_), .CO(
        CARRYB_9__12_), .S(SUMB_9__12_) );
  FA_X1 S2_9_13 ( .A(ab_9__13_), .B(CARRYB_8__13_), .CI(SUMB_8__14_), .CO(
        CARRYB_9__13_), .S(SUMB_9__13_) );
  FA_X1 S2_9_14 ( .A(ab_9__14_), .B(CARRYB_8__14_), .CI(SUMB_8__15_), .CO(
        CARRYB_9__14_), .S(SUMB_9__14_) );
  FA_X1 S2_9_15 ( .A(ab_9__15_), .B(CARRYB_8__15_), .CI(SUMB_8__16_), .CO(
        CARRYB_9__15_), .S(SUMB_9__15_) );
  FA_X1 S2_9_16 ( .A(ab_9__16_), .B(CARRYB_8__16_), .CI(SUMB_8__17_), .CO(
        CARRYB_9__16_), .S(SUMB_9__16_) );
  FA_X1 S2_9_17 ( .A(ab_9__17_), .B(CARRYB_8__17_), .CI(SUMB_8__18_), .CO(
        CARRYB_9__17_), .S(SUMB_9__17_) );
  FA_X1 S2_9_18 ( .A(ab_9__18_), .B(CARRYB_8__18_), .CI(SUMB_8__19_), .CO(
        CARRYB_9__18_), .S(SUMB_9__18_) );
  FA_X1 S2_9_19 ( .A(ab_9__19_), .B(CARRYB_8__19_), .CI(SUMB_8__20_), .CO(
        CARRYB_9__19_), .S(SUMB_9__19_) );
  FA_X1 S2_9_20 ( .A(ab_9__20_), .B(CARRYB_8__20_), .CI(SUMB_8__21_), .CO(
        CARRYB_9__20_), .S(SUMB_9__20_) );
  FA_X1 S2_9_21 ( .A(ab_9__21_), .B(CARRYB_8__21_), .CI(SUMB_8__22_), .CO(
        CARRYB_9__21_), .S(SUMB_9__21_) );
  FA_X1 S3_9_22 ( .A(ab_9__22_), .B(CARRYB_8__22_), .CI(A[8]), .CO(
        CARRYB_9__22_), .S(SUMB_9__22_) );
  FA_X1 S1_8_0 ( .A(ab_8__0_), .B(CARRYB_7__0_), .CI(SUMB_7__1_), .CO(
        CARRYB_8__0_), .S(A1_6_) );
  FA_X1 S2_8_1 ( .A(ab_8__1_), .B(CARRYB_7__1_), .CI(SUMB_7__2_), .CO(
        CARRYB_8__1_), .S(SUMB_8__1_) );
  FA_X1 S2_8_2 ( .A(ab_8__2_), .B(CARRYB_7__2_), .CI(SUMB_7__3_), .CO(
        CARRYB_8__2_), .S(SUMB_8__2_) );
  FA_X1 S2_8_3 ( .A(ab_8__3_), .B(CARRYB_7__3_), .CI(SUMB_7__4_), .CO(
        CARRYB_8__3_), .S(SUMB_8__3_) );
  FA_X1 S2_8_4 ( .A(ab_8__4_), .B(CARRYB_7__4_), .CI(SUMB_7__5_), .CO(
        CARRYB_8__4_), .S(SUMB_8__4_) );
  FA_X1 S2_8_5 ( .A(ab_8__5_), .B(CARRYB_7__5_), .CI(SUMB_7__6_), .CO(
        CARRYB_8__5_), .S(SUMB_8__5_) );
  FA_X1 S2_8_6 ( .A(ab_8__6_), .B(CARRYB_7__6_), .CI(SUMB_7__7_), .CO(
        CARRYB_8__6_), .S(SUMB_8__6_) );
  FA_X1 S2_8_7 ( .A(ab_8__7_), .B(CARRYB_7__7_), .CI(SUMB_7__8_), .CO(
        CARRYB_8__7_), .S(SUMB_8__7_) );
  FA_X1 S2_8_8 ( .A(ab_8__8_), .B(CARRYB_7__8_), .CI(SUMB_7__9_), .CO(
        CARRYB_8__8_), .S(SUMB_8__8_) );
  FA_X1 S2_8_9 ( .A(ab_8__9_), .B(CARRYB_7__9_), .CI(SUMB_7__10_), .CO(
        CARRYB_8__9_), .S(SUMB_8__9_) );
  FA_X1 S2_8_10 ( .A(ab_8__10_), .B(CARRYB_7__10_), .CI(SUMB_7__11_), .CO(
        CARRYB_8__10_), .S(SUMB_8__10_) );
  FA_X1 S2_8_11 ( .A(ab_8__11_), .B(CARRYB_7__11_), .CI(SUMB_7__12_), .CO(
        CARRYB_8__11_), .S(SUMB_8__11_) );
  FA_X1 S2_8_12 ( .A(ab_8__12_), .B(CARRYB_7__12_), .CI(SUMB_7__13_), .CO(
        CARRYB_8__12_), .S(SUMB_8__12_) );
  FA_X1 S2_8_13 ( .A(ab_8__13_), .B(CARRYB_7__13_), .CI(SUMB_7__14_), .CO(
        CARRYB_8__13_), .S(SUMB_8__13_) );
  FA_X1 S2_8_14 ( .A(ab_8__14_), .B(CARRYB_7__14_), .CI(SUMB_7__15_), .CO(
        CARRYB_8__14_), .S(SUMB_8__14_) );
  FA_X1 S2_8_15 ( .A(ab_8__15_), .B(CARRYB_7__15_), .CI(SUMB_7__16_), .CO(
        CARRYB_8__15_), .S(SUMB_8__15_) );
  FA_X1 S2_8_16 ( .A(ab_8__16_), .B(CARRYB_7__16_), .CI(SUMB_7__17_), .CO(
        CARRYB_8__16_), .S(SUMB_8__16_) );
  FA_X1 S2_8_17 ( .A(ab_8__17_), .B(CARRYB_7__17_), .CI(SUMB_7__18_), .CO(
        CARRYB_8__17_), .S(SUMB_8__17_) );
  FA_X1 S2_8_18 ( .A(ab_8__18_), .B(CARRYB_7__18_), .CI(SUMB_7__19_), .CO(
        CARRYB_8__18_), .S(SUMB_8__18_) );
  FA_X1 S2_8_19 ( .A(ab_8__19_), .B(CARRYB_7__19_), .CI(SUMB_7__20_), .CO(
        CARRYB_8__19_), .S(SUMB_8__19_) );
  FA_X1 S2_8_20 ( .A(ab_8__20_), .B(CARRYB_7__20_), .CI(SUMB_7__21_), .CO(
        CARRYB_8__20_), .S(SUMB_8__20_) );
  FA_X1 S2_8_21 ( .A(ab_8__21_), .B(CARRYB_7__21_), .CI(SUMB_7__22_), .CO(
        CARRYB_8__21_), .S(SUMB_8__21_) );
  FA_X1 S3_8_22 ( .A(ab_8__22_), .B(CARRYB_7__22_), .CI(A[7]), .CO(
        CARRYB_8__22_), .S(SUMB_8__22_) );
  FA_X1 S1_7_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(A1_5_) );
  FA_X1 S2_7_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S2_7_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S2_7_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S2_7_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S2_7_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S2_7_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(SUMB_6__7_), .CO(
        CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S2_7_7 ( .A(ab_7__7_), .B(CARRYB_6__7_), .CI(SUMB_6__8_), .CO(
        CARRYB_7__7_), .S(SUMB_7__7_) );
  FA_X1 S2_7_8 ( .A(ab_7__8_), .B(CARRYB_6__8_), .CI(SUMB_6__9_), .CO(
        CARRYB_7__8_), .S(SUMB_7__8_) );
  FA_X1 S2_7_9 ( .A(ab_7__9_), .B(CARRYB_6__9_), .CI(SUMB_6__10_), .CO(
        CARRYB_7__9_), .S(SUMB_7__9_) );
  FA_X1 S2_7_10 ( .A(ab_7__10_), .B(CARRYB_6__10_), .CI(SUMB_6__11_), .CO(
        CARRYB_7__10_), .S(SUMB_7__10_) );
  FA_X1 S2_7_11 ( .A(ab_7__11_), .B(CARRYB_6__11_), .CI(SUMB_6__12_), .CO(
        CARRYB_7__11_), .S(SUMB_7__11_) );
  FA_X1 S2_7_12 ( .A(ab_7__12_), .B(CARRYB_6__12_), .CI(SUMB_6__13_), .CO(
        CARRYB_7__12_), .S(SUMB_7__12_) );
  FA_X1 S2_7_13 ( .A(ab_7__13_), .B(CARRYB_6__13_), .CI(SUMB_6__14_), .CO(
        CARRYB_7__13_), .S(SUMB_7__13_) );
  FA_X1 S2_7_14 ( .A(ab_7__14_), .B(CARRYB_6__14_), .CI(SUMB_6__15_), .CO(
        CARRYB_7__14_), .S(SUMB_7__14_) );
  FA_X1 S2_7_15 ( .A(ab_7__15_), .B(CARRYB_6__15_), .CI(SUMB_6__16_), .CO(
        CARRYB_7__15_), .S(SUMB_7__15_) );
  FA_X1 S2_7_16 ( .A(ab_7__16_), .B(CARRYB_6__16_), .CI(SUMB_6__17_), .CO(
        CARRYB_7__16_), .S(SUMB_7__16_) );
  FA_X1 S2_7_17 ( .A(ab_7__17_), .B(CARRYB_6__17_), .CI(SUMB_6__18_), .CO(
        CARRYB_7__17_), .S(SUMB_7__17_) );
  FA_X1 S2_7_18 ( .A(ab_7__18_), .B(CARRYB_6__18_), .CI(SUMB_6__19_), .CO(
        CARRYB_7__18_), .S(SUMB_7__18_) );
  FA_X1 S2_7_19 ( .A(ab_7__19_), .B(CARRYB_6__19_), .CI(SUMB_6__20_), .CO(
        CARRYB_7__19_), .S(SUMB_7__19_) );
  FA_X1 S2_7_20 ( .A(ab_7__20_), .B(CARRYB_6__20_), .CI(SUMB_6__21_), .CO(
        CARRYB_7__20_), .S(SUMB_7__20_) );
  FA_X1 S2_7_21 ( .A(ab_7__21_), .B(CARRYB_6__21_), .CI(SUMB_6__22_), .CO(
        CARRYB_7__21_), .S(SUMB_7__21_) );
  FA_X1 S3_7_22 ( .A(ab_7__22_), .B(CARRYB_6__22_), .CI(A[6]), .CO(
        CARRYB_7__22_), .S(SUMB_7__22_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S2_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(SUMB_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S2_6_7 ( .A(ab_6__7_), .B(CARRYB_5__7_), .CI(SUMB_5__8_), .CO(
        CARRYB_6__7_), .S(SUMB_6__7_) );
  FA_X1 S2_6_8 ( .A(ab_6__8_), .B(CARRYB_5__8_), .CI(SUMB_5__9_), .CO(
        CARRYB_6__8_), .S(SUMB_6__8_) );
  FA_X1 S2_6_9 ( .A(ab_6__9_), .B(CARRYB_5__9_), .CI(SUMB_5__10_), .CO(
        CARRYB_6__9_), .S(SUMB_6__9_) );
  FA_X1 S2_6_10 ( .A(ab_6__10_), .B(CARRYB_5__10_), .CI(SUMB_5__11_), .CO(
        CARRYB_6__10_), .S(SUMB_6__10_) );
  FA_X1 S2_6_11 ( .A(ab_6__11_), .B(CARRYB_5__11_), .CI(SUMB_5__12_), .CO(
        CARRYB_6__11_), .S(SUMB_6__11_) );
  FA_X1 S2_6_12 ( .A(ab_6__12_), .B(CARRYB_5__12_), .CI(SUMB_5__13_), .CO(
        CARRYB_6__12_), .S(SUMB_6__12_) );
  FA_X1 S2_6_13 ( .A(ab_6__13_), .B(CARRYB_5__13_), .CI(SUMB_5__14_), .CO(
        CARRYB_6__13_), .S(SUMB_6__13_) );
  FA_X1 S2_6_14 ( .A(ab_6__14_), .B(CARRYB_5__14_), .CI(SUMB_5__15_), .CO(
        CARRYB_6__14_), .S(SUMB_6__14_) );
  FA_X1 S2_6_15 ( .A(ab_6__15_), .B(CARRYB_5__15_), .CI(SUMB_5__16_), .CO(
        CARRYB_6__15_), .S(SUMB_6__15_) );
  FA_X1 S2_6_16 ( .A(ab_6__16_), .B(CARRYB_5__16_), .CI(SUMB_5__17_), .CO(
        CARRYB_6__16_), .S(SUMB_6__16_) );
  FA_X1 S2_6_17 ( .A(ab_6__17_), .B(CARRYB_5__17_), .CI(SUMB_5__18_), .CO(
        CARRYB_6__17_), .S(SUMB_6__17_) );
  FA_X1 S2_6_18 ( .A(ab_6__18_), .B(CARRYB_5__18_), .CI(SUMB_5__19_), .CO(
        CARRYB_6__18_), .S(SUMB_6__18_) );
  FA_X1 S2_6_19 ( .A(ab_6__19_), .B(CARRYB_5__19_), .CI(SUMB_5__20_), .CO(
        CARRYB_6__19_), .S(SUMB_6__19_) );
  FA_X1 S2_6_20 ( .A(ab_6__20_), .B(CARRYB_5__20_), .CI(SUMB_5__21_), .CO(
        CARRYB_6__20_), .S(SUMB_6__20_) );
  FA_X1 S2_6_21 ( .A(ab_6__21_), .B(CARRYB_5__21_), .CI(SUMB_5__22_), .CO(
        CARRYB_6__21_), .S(SUMB_6__21_) );
  FA_X1 S3_6_22 ( .A(ab_6__22_), .B(CARRYB_5__22_), .CI(A[5]), .CO(
        CARRYB_6__22_), .S(SUMB_6__22_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S2_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(SUMB_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S2_5_7 ( .A(ab_5__7_), .B(CARRYB_4__7_), .CI(SUMB_4__8_), .CO(
        CARRYB_5__7_), .S(SUMB_5__7_) );
  FA_X1 S2_5_8 ( .A(ab_5__8_), .B(CARRYB_4__8_), .CI(SUMB_4__9_), .CO(
        CARRYB_5__8_), .S(SUMB_5__8_) );
  FA_X1 S2_5_9 ( .A(ab_5__9_), .B(CARRYB_4__9_), .CI(SUMB_4__10_), .CO(
        CARRYB_5__9_), .S(SUMB_5__9_) );
  FA_X1 S2_5_10 ( .A(ab_5__10_), .B(CARRYB_4__10_), .CI(SUMB_4__11_), .CO(
        CARRYB_5__10_), .S(SUMB_5__10_) );
  FA_X1 S2_5_11 ( .A(ab_5__11_), .B(CARRYB_4__11_), .CI(SUMB_4__12_), .CO(
        CARRYB_5__11_), .S(SUMB_5__11_) );
  FA_X1 S2_5_12 ( .A(ab_5__12_), .B(CARRYB_4__12_), .CI(SUMB_4__13_), .CO(
        CARRYB_5__12_), .S(SUMB_5__12_) );
  FA_X1 S2_5_13 ( .A(ab_5__13_), .B(CARRYB_4__13_), .CI(SUMB_4__14_), .CO(
        CARRYB_5__13_), .S(SUMB_5__13_) );
  FA_X1 S2_5_14 ( .A(ab_5__14_), .B(CARRYB_4__14_), .CI(SUMB_4__15_), .CO(
        CARRYB_5__14_), .S(SUMB_5__14_) );
  FA_X1 S2_5_15 ( .A(ab_5__15_), .B(CARRYB_4__15_), .CI(SUMB_4__16_), .CO(
        CARRYB_5__15_), .S(SUMB_5__15_) );
  FA_X1 S2_5_16 ( .A(ab_5__16_), .B(CARRYB_4__16_), .CI(SUMB_4__17_), .CO(
        CARRYB_5__16_), .S(SUMB_5__16_) );
  FA_X1 S2_5_17 ( .A(ab_5__17_), .B(CARRYB_4__17_), .CI(SUMB_4__18_), .CO(
        CARRYB_5__17_), .S(SUMB_5__17_) );
  FA_X1 S2_5_18 ( .A(ab_5__18_), .B(CARRYB_4__18_), .CI(SUMB_4__19_), .CO(
        CARRYB_5__18_), .S(SUMB_5__18_) );
  FA_X1 S2_5_19 ( .A(ab_5__19_), .B(CARRYB_4__19_), .CI(SUMB_4__20_), .CO(
        CARRYB_5__19_), .S(SUMB_5__19_) );
  FA_X1 S2_5_20 ( .A(ab_5__20_), .B(CARRYB_4__20_), .CI(SUMB_4__21_), .CO(
        CARRYB_5__20_), .S(SUMB_5__20_) );
  FA_X1 S2_5_21 ( .A(ab_5__21_), .B(CARRYB_4__21_), .CI(SUMB_4__22_), .CO(
        CARRYB_5__21_), .S(SUMB_5__21_) );
  FA_X1 S3_5_22 ( .A(ab_5__22_), .B(CARRYB_4__22_), .CI(A[4]), .CO(
        CARRYB_5__22_), .S(SUMB_5__22_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S2_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(SUMB_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S2_4_7 ( .A(ab_4__7_), .B(CARRYB_3__7_), .CI(SUMB_3__8_), .CO(
        CARRYB_4__7_), .S(SUMB_4__7_) );
  FA_X1 S2_4_8 ( .A(ab_4__8_), .B(CARRYB_3__8_), .CI(SUMB_3__9_), .CO(
        CARRYB_4__8_), .S(SUMB_4__8_) );
  FA_X1 S2_4_9 ( .A(ab_4__9_), .B(CARRYB_3__9_), .CI(SUMB_3__10_), .CO(
        CARRYB_4__9_), .S(SUMB_4__9_) );
  FA_X1 S2_4_10 ( .A(ab_4__10_), .B(CARRYB_3__10_), .CI(SUMB_3__11_), .CO(
        CARRYB_4__10_), .S(SUMB_4__10_) );
  FA_X1 S2_4_11 ( .A(ab_4__11_), .B(CARRYB_3__11_), .CI(SUMB_3__12_), .CO(
        CARRYB_4__11_), .S(SUMB_4__11_) );
  FA_X1 S2_4_12 ( .A(ab_4__12_), .B(CARRYB_3__12_), .CI(SUMB_3__13_), .CO(
        CARRYB_4__12_), .S(SUMB_4__12_) );
  FA_X1 S2_4_13 ( .A(ab_4__13_), .B(CARRYB_3__13_), .CI(SUMB_3__14_), .CO(
        CARRYB_4__13_), .S(SUMB_4__13_) );
  FA_X1 S2_4_14 ( .A(ab_4__14_), .B(CARRYB_3__14_), .CI(SUMB_3__15_), .CO(
        CARRYB_4__14_), .S(SUMB_4__14_) );
  FA_X1 S2_4_15 ( .A(ab_4__15_), .B(CARRYB_3__15_), .CI(SUMB_3__16_), .CO(
        CARRYB_4__15_), .S(SUMB_4__15_) );
  FA_X1 S2_4_16 ( .A(ab_4__16_), .B(CARRYB_3__16_), .CI(SUMB_3__17_), .CO(
        CARRYB_4__16_), .S(SUMB_4__16_) );
  FA_X1 S2_4_17 ( .A(ab_4__17_), .B(CARRYB_3__17_), .CI(SUMB_3__18_), .CO(
        CARRYB_4__17_), .S(SUMB_4__17_) );
  FA_X1 S2_4_18 ( .A(ab_4__18_), .B(CARRYB_3__18_), .CI(SUMB_3__19_), .CO(
        CARRYB_4__18_), .S(SUMB_4__18_) );
  FA_X1 S2_4_19 ( .A(ab_4__19_), .B(CARRYB_3__19_), .CI(SUMB_3__20_), .CO(
        CARRYB_4__19_), .S(SUMB_4__19_) );
  FA_X1 S2_4_20 ( .A(ab_4__20_), .B(CARRYB_3__20_), .CI(SUMB_3__21_), .CO(
        CARRYB_4__20_), .S(SUMB_4__20_) );
  FA_X1 S2_4_21 ( .A(ab_4__21_), .B(CARRYB_3__21_), .CI(SUMB_3__22_), .CO(
        CARRYB_4__21_), .S(SUMB_4__21_) );
  FA_X1 S3_4_22 ( .A(ab_4__22_), .B(CARRYB_3__22_), .CI(A[3]), .CO(
        CARRYB_4__22_), .S(SUMB_4__22_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S2_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(SUMB_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S2_3_7 ( .A(ab_3__7_), .B(CARRYB_2__7_), .CI(SUMB_2__8_), .CO(
        CARRYB_3__7_), .S(SUMB_3__7_) );
  FA_X1 S2_3_8 ( .A(ab_3__8_), .B(CARRYB_2__8_), .CI(SUMB_2__9_), .CO(
        CARRYB_3__8_), .S(SUMB_3__8_) );
  FA_X1 S2_3_9 ( .A(ab_3__9_), .B(CARRYB_2__9_), .CI(SUMB_2__10_), .CO(
        CARRYB_3__9_), .S(SUMB_3__9_) );
  FA_X1 S2_3_10 ( .A(ab_3__10_), .B(CARRYB_2__10_), .CI(SUMB_2__11_), .CO(
        CARRYB_3__10_), .S(SUMB_3__10_) );
  FA_X1 S2_3_11 ( .A(ab_3__11_), .B(CARRYB_2__11_), .CI(SUMB_2__12_), .CO(
        CARRYB_3__11_), .S(SUMB_3__11_) );
  FA_X1 S2_3_12 ( .A(ab_3__12_), .B(CARRYB_2__12_), .CI(SUMB_2__13_), .CO(
        CARRYB_3__12_), .S(SUMB_3__12_) );
  FA_X1 S2_3_13 ( .A(ab_3__13_), .B(CARRYB_2__13_), .CI(SUMB_2__14_), .CO(
        CARRYB_3__13_), .S(SUMB_3__13_) );
  FA_X1 S2_3_14 ( .A(ab_3__14_), .B(CARRYB_2__14_), .CI(SUMB_2__15_), .CO(
        CARRYB_3__14_), .S(SUMB_3__14_) );
  FA_X1 S2_3_15 ( .A(ab_3__15_), .B(CARRYB_2__15_), .CI(SUMB_2__16_), .CO(
        CARRYB_3__15_), .S(SUMB_3__15_) );
  FA_X1 S2_3_16 ( .A(ab_3__16_), .B(CARRYB_2__16_), .CI(SUMB_2__17_), .CO(
        CARRYB_3__16_), .S(SUMB_3__16_) );
  FA_X1 S2_3_17 ( .A(ab_3__17_), .B(CARRYB_2__17_), .CI(SUMB_2__18_), .CO(
        CARRYB_3__17_), .S(SUMB_3__17_) );
  FA_X1 S2_3_18 ( .A(ab_3__18_), .B(CARRYB_2__18_), .CI(SUMB_2__19_), .CO(
        CARRYB_3__18_), .S(SUMB_3__18_) );
  FA_X1 S2_3_19 ( .A(ab_3__19_), .B(CARRYB_2__19_), .CI(SUMB_2__20_), .CO(
        CARRYB_3__19_), .S(SUMB_3__19_) );
  FA_X1 S2_3_20 ( .A(ab_3__20_), .B(CARRYB_2__20_), .CI(SUMB_2__21_), .CO(
        CARRYB_3__20_), .S(SUMB_3__20_) );
  FA_X1 S2_3_21 ( .A(ab_3__21_), .B(CARRYB_2__21_), .CI(SUMB_2__22_), .CO(
        CARRYB_3__21_), .S(SUMB_3__21_) );
  FA_X1 S3_3_22 ( .A(ab_3__22_), .B(CARRYB_2__22_), .CI(A[2]), .CO(
        CARRYB_3__22_), .S(SUMB_3__22_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(CARRYB_1__0_), .CI(n26), .CO(CARRYB_2__0_), 
        .S(A1_0_) );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n5), .CI(n25), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n4), .CI(n24), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n3), .CI(n23), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n2), .CI(n27), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n16), .CI(n37), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S2_2_6 ( .A(ab_2__6_), .B(n15), .CI(n36), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  FA_X1 S2_2_7 ( .A(ab_2__7_), .B(n14), .CI(n35), .CO(CARRYB_2__7_), .S(
        SUMB_2__7_) );
  FA_X1 S2_2_8 ( .A(ab_2__8_), .B(n13), .CI(n34), .CO(CARRYB_2__8_), .S(
        SUMB_2__8_) );
  FA_X1 S2_2_9 ( .A(ab_2__9_), .B(n12), .CI(n33), .CO(CARRYB_2__9_), .S(
        SUMB_2__9_) );
  FA_X1 S2_2_10 ( .A(ab_2__10_), .B(n11), .CI(n32), .CO(CARRYB_2__10_), .S(
        SUMB_2__10_) );
  FA_X1 S2_2_11 ( .A(ab_2__11_), .B(n10), .CI(n31), .CO(CARRYB_2__11_), .S(
        SUMB_2__11_) );
  FA_X1 S2_2_12 ( .A(ab_2__12_), .B(n9), .CI(n30), .CO(CARRYB_2__12_), .S(
        SUMB_2__12_) );
  FA_X1 S2_2_13 ( .A(ab_2__13_), .B(n8), .CI(n29), .CO(CARRYB_2__13_), .S(
        SUMB_2__13_) );
  FA_X1 S2_2_14 ( .A(ab_2__14_), .B(n7), .CI(n28), .CO(CARRYB_2__14_), .S(
        SUMB_2__14_) );
  FA_X1 S2_2_15 ( .A(ab_2__15_), .B(n6), .CI(n40), .CO(CARRYB_2__15_), .S(
        SUMB_2__15_) );
  FA_X1 S2_2_16 ( .A(ab_2__16_), .B(n19), .CI(n39), .CO(CARRYB_2__16_), .S(
        SUMB_2__16_) );
  FA_X1 S2_2_17 ( .A(ab_2__17_), .B(n18), .CI(n38), .CO(CARRYB_2__17_), .S(
        SUMB_2__17_) );
  FA_X1 S2_2_18 ( .A(ab_2__18_), .B(n17), .CI(n44), .CO(CARRYB_2__18_), .S(
        SUMB_2__18_) );
  FA_X1 S2_2_19 ( .A(ab_2__19_), .B(n22), .CI(n43), .CO(CARRYB_2__19_), .S(
        SUMB_2__19_) );
  FA_X1 S2_2_20 ( .A(ab_2__20_), .B(n21), .CI(n42), .CO(CARRYB_2__20_), .S(
        SUMB_2__20_) );
  FA_X1 S2_2_21 ( .A(ab_2__21_), .B(n20), .CI(n41), .CO(CARRYB_2__21_), .S(
        SUMB_2__21_) );
  FA_X1 S3_2_22 ( .A(ab_2__22_), .B(n45), .CI(A[1]), .CO(CARRYB_2__22_), .S(
        SUMB_2__22_) );
  FPM_DW01_add_2 FS_1 ( .A({1'b0, n98, n84, n87, n83, n65, n53, n71, n52, n67, 
        n51, n70, n50, n69, n49, n66, n48, n68, n47, n63, n46, n64, n72, n82, 
        SUMB_23__0_, A1_20_, A1_19_, A1_18_, A1_17_, A1_16_, A1_15_, A1_14_, 
        A1_13_, A1_12_, A1_11_, A1_10_, A1_9_, A1_8_, A1_7_, A1_6_, A1_5_, 
        A1_4_, A1_3_, A1_2_, A1_1_, A1_0_}), .B({CARRYB_23__22_, n89, n86, n88, 
        n85, n75, n62, n81, n61, n77, n60, n80, n59, n79, n58, n76, n57, n78, 
        n56, n73, n55, n74, n54, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({PRODUCT[47:23], 
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21}) );
  AND2_X1 U2 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n2) );
  AND2_X1 U3 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n3) );
  AND2_X1 U4 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n4) );
  AND2_X1 U5 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n5) );
  AND2_X1 U6 ( .A1(ab_0__16_), .A2(ab_1__15_), .ZN(n6) );
  AND2_X1 U7 ( .A1(ab_0__15_), .A2(ab_1__14_), .ZN(n7) );
  AND2_X1 U8 ( .A1(ab_0__14_), .A2(ab_1__13_), .ZN(n8) );
  AND2_X1 U9 ( .A1(ab_0__13_), .A2(ab_1__12_), .ZN(n9) );
  AND2_X1 U10 ( .A1(ab_0__12_), .A2(ab_1__11_), .ZN(n10) );
  AND2_X1 U11 ( .A1(ab_0__11_), .A2(ab_1__10_), .ZN(n11) );
  AND2_X1 U12 ( .A1(ab_0__10_), .A2(ab_1__9_), .ZN(n12) );
  AND2_X1 U13 ( .A1(ab_0__9_), .A2(ab_1__8_), .ZN(n13) );
  AND2_X1 U14 ( .A1(ab_0__8_), .A2(ab_1__7_), .ZN(n14) );
  AND2_X1 U15 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n15) );
  AND2_X1 U16 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n16) );
  AND2_X1 U17 ( .A1(ab_0__19_), .A2(ab_1__18_), .ZN(n17) );
  AND2_X1 U18 ( .A1(ab_0__18_), .A2(ab_1__17_), .ZN(n18) );
  AND2_X1 U19 ( .A1(ab_0__17_), .A2(ab_1__16_), .ZN(n19) );
  AND2_X1 U20 ( .A1(ab_0__22_), .A2(ab_1__21_), .ZN(n20) );
  AND2_X1 U21 ( .A1(ab_0__21_), .A2(ab_1__20_), .ZN(n21) );
  AND2_X1 U22 ( .A1(ab_0__20_), .A2(ab_1__19_), .ZN(n22) );
  XOR2_X1 U23 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n23) );
  XOR2_X1 U24 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n24) );
  XOR2_X1 U25 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n25) );
  XOR2_X1 U26 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n26) );
  XOR2_X1 U27 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n27) );
  XOR2_X1 U28 ( .A(ab_1__15_), .B(ab_0__16_), .Z(n28) );
  XOR2_X1 U29 ( .A(ab_1__14_), .B(ab_0__15_), .Z(n29) );
  XOR2_X1 U30 ( .A(ab_1__13_), .B(ab_0__14_), .Z(n30) );
  XOR2_X1 U31 ( .A(ab_1__12_), .B(ab_0__13_), .Z(n31) );
  XOR2_X1 U32 ( .A(ab_1__11_), .B(ab_0__12_), .Z(n32) );
  XOR2_X1 U33 ( .A(ab_1__10_), .B(ab_0__11_), .Z(n33) );
  XOR2_X1 U34 ( .A(ab_1__9_), .B(ab_0__10_), .Z(n34) );
  XOR2_X1 U35 ( .A(ab_1__8_), .B(ab_0__9_), .Z(n35) );
  XOR2_X1 U36 ( .A(ab_1__7_), .B(ab_0__8_), .Z(n36) );
  XOR2_X1 U37 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n37) );
  XOR2_X1 U38 ( .A(ab_1__18_), .B(ab_0__19_), .Z(n38) );
  XOR2_X1 U39 ( .A(ab_1__17_), .B(ab_0__18_), .Z(n39) );
  XOR2_X1 U40 ( .A(ab_1__16_), .B(ab_0__17_), .Z(n40) );
  XOR2_X1 U41 ( .A(ab_1__22_), .B(n95), .Z(n41) );
  XOR2_X1 U42 ( .A(ab_1__21_), .B(ab_0__22_), .Z(n42) );
  XOR2_X1 U43 ( .A(ab_1__20_), .B(ab_0__21_), .Z(n43) );
  XOR2_X1 U44 ( .A(ab_1__19_), .B(ab_0__20_), .Z(n44) );
  AND2_X1 U45 ( .A1(n95), .A2(ab_1__22_), .ZN(n45) );
  XOR2_X1 U46 ( .A(CARRYB_23__3_), .B(SUMB_23__4_), .Z(n46) );
  XOR2_X1 U47 ( .A(CARRYB_23__5_), .B(SUMB_23__6_), .Z(n47) );
  XOR2_X1 U48 ( .A(CARRYB_23__7_), .B(SUMB_23__8_), .Z(n48) );
  XOR2_X1 U49 ( .A(CARRYB_23__9_), .B(SUMB_23__10_), .Z(n49) );
  XOR2_X1 U50 ( .A(CARRYB_23__11_), .B(SUMB_23__12_), .Z(n50) );
  XOR2_X1 U51 ( .A(CARRYB_23__13_), .B(SUMB_23__14_), .Z(n51) );
  XOR2_X1 U52 ( .A(CARRYB_23__15_), .B(SUMB_23__16_), .Z(n52) );
  XOR2_X1 U53 ( .A(CARRYB_23__17_), .B(SUMB_23__18_), .Z(n53) );
  AND2_X1 U54 ( .A1(CARRYB_23__0_), .A2(SUMB_23__1_), .ZN(n54) );
  AND2_X1 U55 ( .A1(CARRYB_23__2_), .A2(SUMB_23__3_), .ZN(n55) );
  AND2_X1 U56 ( .A1(CARRYB_23__4_), .A2(SUMB_23__5_), .ZN(n56) );
  AND2_X1 U57 ( .A1(CARRYB_23__6_), .A2(SUMB_23__7_), .ZN(n57) );
  AND2_X1 U58 ( .A1(CARRYB_23__8_), .A2(SUMB_23__9_), .ZN(n58) );
  AND2_X1 U59 ( .A1(CARRYB_23__10_), .A2(SUMB_23__11_), .ZN(n59) );
  AND2_X1 U60 ( .A1(CARRYB_23__12_), .A2(SUMB_23__13_), .ZN(n60) );
  AND2_X1 U61 ( .A1(CARRYB_23__14_), .A2(SUMB_23__15_), .ZN(n61) );
  AND2_X1 U62 ( .A1(CARRYB_23__16_), .A2(SUMB_23__17_), .ZN(n62) );
  XOR2_X1 U63 ( .A(CARRYB_23__4_), .B(SUMB_23__5_), .Z(n63) );
  XOR2_X1 U64 ( .A(CARRYB_23__2_), .B(SUMB_23__3_), .Z(n64) );
  XOR2_X1 U65 ( .A(CARRYB_23__18_), .B(SUMB_23__19_), .Z(n65) );
  XOR2_X1 U66 ( .A(CARRYB_23__8_), .B(SUMB_23__9_), .Z(n66) );
  XOR2_X1 U67 ( .A(CARRYB_23__14_), .B(SUMB_23__15_), .Z(n67) );
  XOR2_X1 U68 ( .A(CARRYB_23__6_), .B(SUMB_23__7_), .Z(n68) );
  XOR2_X1 U69 ( .A(CARRYB_23__10_), .B(SUMB_23__11_), .Z(n69) );
  XOR2_X1 U70 ( .A(CARRYB_23__12_), .B(SUMB_23__13_), .Z(n70) );
  XOR2_X1 U71 ( .A(CARRYB_23__16_), .B(SUMB_23__17_), .Z(n71) );
  XOR2_X1 U72 ( .A(CARRYB_23__1_), .B(SUMB_23__2_), .Z(n72) );
  AND2_X1 U73 ( .A1(CARRYB_23__3_), .A2(SUMB_23__4_), .ZN(n73) );
  AND2_X1 U74 ( .A1(CARRYB_23__1_), .A2(SUMB_23__2_), .ZN(n74) );
  AND2_X1 U75 ( .A1(CARRYB_23__17_), .A2(SUMB_23__18_), .ZN(n75) );
  AND2_X1 U76 ( .A1(CARRYB_23__7_), .A2(SUMB_23__8_), .ZN(n76) );
  AND2_X1 U77 ( .A1(CARRYB_23__13_), .A2(SUMB_23__14_), .ZN(n77) );
  AND2_X1 U78 ( .A1(CARRYB_23__5_), .A2(SUMB_23__6_), .ZN(n78) );
  AND2_X1 U79 ( .A1(CARRYB_23__9_), .A2(SUMB_23__10_), .ZN(n79) );
  AND2_X1 U80 ( .A1(CARRYB_23__11_), .A2(SUMB_23__12_), .ZN(n80) );
  AND2_X1 U81 ( .A1(CARRYB_23__15_), .A2(SUMB_23__16_), .ZN(n81) );
  XOR2_X1 U82 ( .A(CARRYB_23__0_), .B(SUMB_23__1_), .Z(n82) );
  INV_X1 U83 ( .A(CARRYB_23__22_), .ZN(n98) );
  XOR2_X1 U84 ( .A(CARRYB_23__19_), .B(SUMB_23__20_), .Z(n83) );
  XOR2_X1 U85 ( .A(CARRYB_23__21_), .B(SUMB_23__22_), .Z(n84) );
  AND2_X1 U86 ( .A1(CARRYB_23__18_), .A2(SUMB_23__19_), .ZN(n85) );
  AND2_X1 U87 ( .A1(CARRYB_23__20_), .A2(SUMB_23__21_), .ZN(n86) );
  XOR2_X1 U88 ( .A(CARRYB_23__20_), .B(SUMB_23__21_), .Z(n87) );
  AND2_X1 U89 ( .A1(CARRYB_23__19_), .A2(SUMB_23__20_), .ZN(n88) );
  AND2_X1 U90 ( .A1(CARRYB_23__21_), .A2(SUMB_23__22_), .ZN(n89) );
  INV_X1 U91 ( .A(A[9]), .ZN(n133) );
  INV_X1 U92 ( .A(B[2]), .ZN(n117) );
  INV_X1 U93 ( .A(B[5]), .ZN(n114) );
  INV_X1 U94 ( .A(B[4]), .ZN(n115) );
  INV_X1 U95 ( .A(B[3]), .ZN(n116) );
  INV_X1 U96 ( .A(A[4]), .ZN(n138) );
  INV_X1 U97 ( .A(A[6]), .ZN(n136) );
  INV_X1 U98 ( .A(A[5]), .ZN(n137) );
  INV_X1 U99 ( .A(A[8]), .ZN(n134) );
  INV_X1 U100 ( .A(A[7]), .ZN(n135) );
  INV_X1 U101 ( .A(A[10]), .ZN(n132) );
  INV_X1 U102 ( .A(B[1]), .ZN(n118) );
  INV_X1 U103 ( .A(B[0]), .ZN(n119) );
  INV_X1 U104 ( .A(A[12]), .ZN(n130) );
  INV_X1 U105 ( .A(A[14]), .ZN(n128) );
  INV_X1 U106 ( .A(A[13]), .ZN(n129) );
  INV_X1 U107 ( .A(A[16]), .ZN(n126) );
  INV_X1 U108 ( .A(A[15]), .ZN(n127) );
  INV_X1 U109 ( .A(A[18]), .ZN(n124) );
  INV_X1 U110 ( .A(A[17]), .ZN(n125) );
  INV_X1 U111 ( .A(A[19]), .ZN(n123) );
  INV_X1 U112 ( .A(A[11]), .ZN(n131) );
  INV_X1 U113 ( .A(A[20]), .ZN(n122) );
  INV_X1 U114 ( .A(A[21]), .ZN(n121) );
  INV_X1 U115 ( .A(A[22]), .ZN(n120) );
  BUF_X4 U116 ( .A(n101), .Z(n90) );
  INV_X1 U117 ( .A(B[19]), .ZN(n101) );
  CLKBUF_X1 U118 ( .A(n102), .Z(n91) );
  BUF_X4 U119 ( .A(n102), .Z(n92) );
  INV_X1 U120 ( .A(B[17]), .ZN(n102) );
  CLKBUF_X1 U121 ( .A(n141), .Z(n93) );
  INV_X1 U122 ( .A(A[0]), .ZN(n141) );
  INV_X2 U123 ( .A(B[18]), .ZN(n94) );
  CLKBUF_X1 U124 ( .A(A[0]), .Z(n95) );
  AND2_X1 U125 ( .A1(B[21]), .A2(A[1]), .ZN(ab_1__21_) );
  AND2_X1 U126 ( .A1(B[20]), .A2(A[0]), .ZN(ab_0__20_) );
  AND2_X1 U127 ( .A1(B[19]), .A2(A[1]), .ZN(ab_1__19_) );
  AND2_X1 U128 ( .A1(B[20]), .A2(A[1]), .ZN(ab_1__20_) );
  AND2_X1 U129 ( .A1(B[21]), .A2(A[0]), .ZN(ab_0__21_) );
  INV_X2 U130 ( .A(B[21]), .ZN(n96) );
  AND2_X1 U131 ( .A1(B[22]), .A2(A[0]), .ZN(ab_0__22_) );
  INV_X1 U132 ( .A(B[22]), .ZN(n99) );
  INV_X1 U133 ( .A(A[1]), .ZN(n97) );
  INV_X2 U134 ( .A(B[20]), .ZN(n100) );
  INV_X2 U135 ( .A(B[16]), .ZN(n103) );
  INV_X2 U136 ( .A(B[15]), .ZN(n104) );
  INV_X2 U137 ( .A(B[14]), .ZN(n105) );
  INV_X2 U138 ( .A(B[13]), .ZN(n106) );
  INV_X2 U139 ( .A(B[12]), .ZN(n107) );
  INV_X2 U140 ( .A(B[11]), .ZN(n108) );
  INV_X2 U141 ( .A(B[10]), .ZN(n109) );
  INV_X2 U142 ( .A(B[9]), .ZN(n110) );
  INV_X2 U143 ( .A(B[8]), .ZN(n111) );
  INV_X2 U144 ( .A(B[7]), .ZN(n112) );
  INV_X2 U145 ( .A(B[6]), .ZN(n113) );
  INV_X2 U146 ( .A(A[3]), .ZN(n139) );
  INV_X2 U147 ( .A(A[2]), .ZN(n140) );
  NOR2_X1 U149 ( .A1(n133), .A2(n110), .ZN(ab_9__9_) );
  NOR2_X1 U150 ( .A1(n133), .A2(n111), .ZN(ab_9__8_) );
  NOR2_X1 U151 ( .A1(n133), .A2(n112), .ZN(ab_9__7_) );
  NOR2_X1 U152 ( .A1(n133), .A2(n113), .ZN(ab_9__6_) );
  NOR2_X1 U153 ( .A1(n133), .A2(n114), .ZN(ab_9__5_) );
  NOR2_X1 U154 ( .A1(n133), .A2(n115), .ZN(ab_9__4_) );
  NOR2_X1 U155 ( .A1(n133), .A2(n116), .ZN(ab_9__3_) );
  NOR2_X1 U156 ( .A1(n133), .A2(n117), .ZN(ab_9__2_) );
  NOR2_X1 U157 ( .A1(n133), .A2(n99), .ZN(ab_9__22_) );
  NOR2_X1 U158 ( .A1(n133), .A2(n96), .ZN(ab_9__21_) );
  NOR2_X1 U159 ( .A1(n133), .A2(n100), .ZN(ab_9__20_) );
  NOR2_X1 U160 ( .A1(n133), .A2(n118), .ZN(ab_9__1_) );
  NOR2_X1 U161 ( .A1(n133), .A2(n90), .ZN(ab_9__19_) );
  NOR2_X1 U162 ( .A1(n133), .A2(n94), .ZN(ab_9__18_) );
  NOR2_X1 U163 ( .A1(n133), .A2(n92), .ZN(ab_9__17_) );
  NOR2_X1 U164 ( .A1(n133), .A2(n103), .ZN(ab_9__16_) );
  NOR2_X1 U165 ( .A1(n133), .A2(n104), .ZN(ab_9__15_) );
  NOR2_X1 U166 ( .A1(n133), .A2(n105), .ZN(ab_9__14_) );
  NOR2_X1 U167 ( .A1(n133), .A2(n106), .ZN(ab_9__13_) );
  NOR2_X1 U168 ( .A1(n133), .A2(n107), .ZN(ab_9__12_) );
  NOR2_X1 U169 ( .A1(n133), .A2(n108), .ZN(ab_9__11_) );
  NOR2_X1 U170 ( .A1(n133), .A2(n109), .ZN(ab_9__10_) );
  NOR2_X1 U171 ( .A1(n133), .A2(n119), .ZN(ab_9__0_) );
  NOR2_X1 U172 ( .A1(n110), .A2(n134), .ZN(ab_8__9_) );
  NOR2_X1 U173 ( .A1(n111), .A2(n134), .ZN(ab_8__8_) );
  NOR2_X1 U174 ( .A1(n112), .A2(n134), .ZN(ab_8__7_) );
  NOR2_X1 U175 ( .A1(n113), .A2(n134), .ZN(ab_8__6_) );
  NOR2_X1 U176 ( .A1(n114), .A2(n134), .ZN(ab_8__5_) );
  NOR2_X1 U177 ( .A1(n115), .A2(n134), .ZN(ab_8__4_) );
  NOR2_X1 U178 ( .A1(n116), .A2(n134), .ZN(ab_8__3_) );
  NOR2_X1 U179 ( .A1(n117), .A2(n134), .ZN(ab_8__2_) );
  NOR2_X1 U180 ( .A1(n99), .A2(n134), .ZN(ab_8__22_) );
  NOR2_X1 U181 ( .A1(n96), .A2(n134), .ZN(ab_8__21_) );
  NOR2_X1 U182 ( .A1(n100), .A2(n134), .ZN(ab_8__20_) );
  NOR2_X1 U183 ( .A1(n118), .A2(n134), .ZN(ab_8__1_) );
  NOR2_X1 U184 ( .A1(n90), .A2(n134), .ZN(ab_8__19_) );
  NOR2_X1 U185 ( .A1(n94), .A2(n134), .ZN(ab_8__18_) );
  NOR2_X1 U186 ( .A1(n92), .A2(n134), .ZN(ab_8__17_) );
  NOR2_X1 U187 ( .A1(n103), .A2(n134), .ZN(ab_8__16_) );
  NOR2_X1 U188 ( .A1(n104), .A2(n134), .ZN(ab_8__15_) );
  NOR2_X1 U189 ( .A1(n105), .A2(n134), .ZN(ab_8__14_) );
  NOR2_X1 U190 ( .A1(n106), .A2(n134), .ZN(ab_8__13_) );
  NOR2_X1 U191 ( .A1(n107), .A2(n134), .ZN(ab_8__12_) );
  NOR2_X1 U192 ( .A1(n108), .A2(n134), .ZN(ab_8__11_) );
  NOR2_X1 U193 ( .A1(n109), .A2(n134), .ZN(ab_8__10_) );
  NOR2_X1 U194 ( .A1(n119), .A2(n134), .ZN(ab_8__0_) );
  NOR2_X1 U195 ( .A1(n110), .A2(n135), .ZN(ab_7__9_) );
  NOR2_X1 U196 ( .A1(n111), .A2(n135), .ZN(ab_7__8_) );
  NOR2_X1 U197 ( .A1(n112), .A2(n135), .ZN(ab_7__7_) );
  NOR2_X1 U198 ( .A1(n113), .A2(n135), .ZN(ab_7__6_) );
  NOR2_X1 U199 ( .A1(n114), .A2(n135), .ZN(ab_7__5_) );
  NOR2_X1 U200 ( .A1(n115), .A2(n135), .ZN(ab_7__4_) );
  NOR2_X1 U201 ( .A1(n116), .A2(n135), .ZN(ab_7__3_) );
  NOR2_X1 U202 ( .A1(n117), .A2(n135), .ZN(ab_7__2_) );
  NOR2_X1 U203 ( .A1(n99), .A2(n135), .ZN(ab_7__22_) );
  NOR2_X1 U204 ( .A1(n96), .A2(n135), .ZN(ab_7__21_) );
  NOR2_X1 U205 ( .A1(n100), .A2(n135), .ZN(ab_7__20_) );
  NOR2_X1 U206 ( .A1(n118), .A2(n135), .ZN(ab_7__1_) );
  NOR2_X1 U207 ( .A1(n90), .A2(n135), .ZN(ab_7__19_) );
  NOR2_X1 U208 ( .A1(n94), .A2(n135), .ZN(ab_7__18_) );
  NOR2_X1 U209 ( .A1(n92), .A2(n135), .ZN(ab_7__17_) );
  NOR2_X1 U210 ( .A1(n103), .A2(n135), .ZN(ab_7__16_) );
  NOR2_X1 U211 ( .A1(n104), .A2(n135), .ZN(ab_7__15_) );
  NOR2_X1 U212 ( .A1(n105), .A2(n135), .ZN(ab_7__14_) );
  NOR2_X1 U213 ( .A1(n106), .A2(n135), .ZN(ab_7__13_) );
  NOR2_X1 U214 ( .A1(n107), .A2(n135), .ZN(ab_7__12_) );
  NOR2_X1 U215 ( .A1(n108), .A2(n135), .ZN(ab_7__11_) );
  NOR2_X1 U216 ( .A1(n109), .A2(n135), .ZN(ab_7__10_) );
  NOR2_X1 U217 ( .A1(n119), .A2(n135), .ZN(ab_7__0_) );
  NOR2_X1 U218 ( .A1(n110), .A2(n136), .ZN(ab_6__9_) );
  NOR2_X1 U219 ( .A1(n111), .A2(n136), .ZN(ab_6__8_) );
  NOR2_X1 U220 ( .A1(n112), .A2(n136), .ZN(ab_6__7_) );
  NOR2_X1 U221 ( .A1(n113), .A2(n136), .ZN(ab_6__6_) );
  NOR2_X1 U222 ( .A1(n114), .A2(n136), .ZN(ab_6__5_) );
  NOR2_X1 U223 ( .A1(n115), .A2(n136), .ZN(ab_6__4_) );
  NOR2_X1 U224 ( .A1(n116), .A2(n136), .ZN(ab_6__3_) );
  NOR2_X1 U225 ( .A1(n117), .A2(n136), .ZN(ab_6__2_) );
  NOR2_X1 U226 ( .A1(n99), .A2(n136), .ZN(ab_6__22_) );
  NOR2_X1 U227 ( .A1(n96), .A2(n136), .ZN(ab_6__21_) );
  NOR2_X1 U228 ( .A1(n100), .A2(n136), .ZN(ab_6__20_) );
  NOR2_X1 U229 ( .A1(n118), .A2(n136), .ZN(ab_6__1_) );
  NOR2_X1 U230 ( .A1(n90), .A2(n136), .ZN(ab_6__19_) );
  NOR2_X1 U231 ( .A1(n94), .A2(n136), .ZN(ab_6__18_) );
  NOR2_X1 U232 ( .A1(n92), .A2(n136), .ZN(ab_6__17_) );
  NOR2_X1 U233 ( .A1(n103), .A2(n136), .ZN(ab_6__16_) );
  NOR2_X1 U234 ( .A1(n104), .A2(n136), .ZN(ab_6__15_) );
  NOR2_X1 U235 ( .A1(n105), .A2(n136), .ZN(ab_6__14_) );
  NOR2_X1 U236 ( .A1(n106), .A2(n136), .ZN(ab_6__13_) );
  NOR2_X1 U237 ( .A1(n107), .A2(n136), .ZN(ab_6__12_) );
  NOR2_X1 U238 ( .A1(n108), .A2(n136), .ZN(ab_6__11_) );
  NOR2_X1 U239 ( .A1(n109), .A2(n136), .ZN(ab_6__10_) );
  NOR2_X1 U240 ( .A1(n119), .A2(n136), .ZN(ab_6__0_) );
  NOR2_X1 U241 ( .A1(n110), .A2(n137), .ZN(ab_5__9_) );
  NOR2_X1 U242 ( .A1(n111), .A2(n137), .ZN(ab_5__8_) );
  NOR2_X1 U243 ( .A1(n112), .A2(n137), .ZN(ab_5__7_) );
  NOR2_X1 U244 ( .A1(n113), .A2(n137), .ZN(ab_5__6_) );
  NOR2_X1 U245 ( .A1(n114), .A2(n137), .ZN(ab_5__5_) );
  NOR2_X1 U246 ( .A1(n115), .A2(n137), .ZN(ab_5__4_) );
  NOR2_X1 U247 ( .A1(n116), .A2(n137), .ZN(ab_5__3_) );
  NOR2_X1 U248 ( .A1(n117), .A2(n137), .ZN(ab_5__2_) );
  NOR2_X1 U249 ( .A1(n99), .A2(n137), .ZN(ab_5__22_) );
  NOR2_X1 U250 ( .A1(n96), .A2(n137), .ZN(ab_5__21_) );
  NOR2_X1 U251 ( .A1(n100), .A2(n137), .ZN(ab_5__20_) );
  NOR2_X1 U252 ( .A1(n118), .A2(n137), .ZN(ab_5__1_) );
  NOR2_X1 U253 ( .A1(n90), .A2(n137), .ZN(ab_5__19_) );
  NOR2_X1 U254 ( .A1(n94), .A2(n137), .ZN(ab_5__18_) );
  NOR2_X1 U255 ( .A1(n92), .A2(n137), .ZN(ab_5__17_) );
  NOR2_X1 U256 ( .A1(n103), .A2(n137), .ZN(ab_5__16_) );
  NOR2_X1 U257 ( .A1(n104), .A2(n137), .ZN(ab_5__15_) );
  NOR2_X1 U258 ( .A1(n105), .A2(n137), .ZN(ab_5__14_) );
  NOR2_X1 U259 ( .A1(n106), .A2(n137), .ZN(ab_5__13_) );
  NOR2_X1 U260 ( .A1(n107), .A2(n137), .ZN(ab_5__12_) );
  NOR2_X1 U261 ( .A1(n108), .A2(n137), .ZN(ab_5__11_) );
  NOR2_X1 U262 ( .A1(n109), .A2(n137), .ZN(ab_5__10_) );
  NOR2_X1 U263 ( .A1(n119), .A2(n137), .ZN(ab_5__0_) );
  NOR2_X1 U264 ( .A1(n110), .A2(n138), .ZN(ab_4__9_) );
  NOR2_X1 U265 ( .A1(n111), .A2(n138), .ZN(ab_4__8_) );
  NOR2_X1 U266 ( .A1(n112), .A2(n138), .ZN(ab_4__7_) );
  NOR2_X1 U267 ( .A1(n113), .A2(n138), .ZN(ab_4__6_) );
  NOR2_X1 U268 ( .A1(n114), .A2(n138), .ZN(ab_4__5_) );
  NOR2_X1 U269 ( .A1(n115), .A2(n138), .ZN(ab_4__4_) );
  NOR2_X1 U270 ( .A1(n116), .A2(n138), .ZN(ab_4__3_) );
  NOR2_X1 U271 ( .A1(n117), .A2(n138), .ZN(ab_4__2_) );
  NOR2_X1 U272 ( .A1(n99), .A2(n138), .ZN(ab_4__22_) );
  NOR2_X1 U273 ( .A1(n96), .A2(n138), .ZN(ab_4__21_) );
  NOR2_X1 U274 ( .A1(n100), .A2(n138), .ZN(ab_4__20_) );
  NOR2_X1 U275 ( .A1(n118), .A2(n138), .ZN(ab_4__1_) );
  NOR2_X1 U276 ( .A1(n90), .A2(n138), .ZN(ab_4__19_) );
  NOR2_X1 U277 ( .A1(n94), .A2(n138), .ZN(ab_4__18_) );
  NOR2_X1 U278 ( .A1(n92), .A2(n138), .ZN(ab_4__17_) );
  NOR2_X1 U279 ( .A1(n103), .A2(n138), .ZN(ab_4__16_) );
  NOR2_X1 U280 ( .A1(n104), .A2(n138), .ZN(ab_4__15_) );
  NOR2_X1 U281 ( .A1(n105), .A2(n138), .ZN(ab_4__14_) );
  NOR2_X1 U282 ( .A1(n106), .A2(n138), .ZN(ab_4__13_) );
  NOR2_X1 U283 ( .A1(n107), .A2(n138), .ZN(ab_4__12_) );
  NOR2_X1 U284 ( .A1(n108), .A2(n138), .ZN(ab_4__11_) );
  NOR2_X1 U285 ( .A1(n109), .A2(n138), .ZN(ab_4__10_) );
  NOR2_X1 U286 ( .A1(n119), .A2(n138), .ZN(ab_4__0_) );
  NOR2_X1 U287 ( .A1(n110), .A2(n139), .ZN(ab_3__9_) );
  NOR2_X1 U288 ( .A1(n111), .A2(n139), .ZN(ab_3__8_) );
  NOR2_X1 U289 ( .A1(n112), .A2(n139), .ZN(ab_3__7_) );
  NOR2_X1 U290 ( .A1(n113), .A2(n139), .ZN(ab_3__6_) );
  NOR2_X1 U291 ( .A1(n114), .A2(n139), .ZN(ab_3__5_) );
  NOR2_X1 U292 ( .A1(n115), .A2(n139), .ZN(ab_3__4_) );
  NOR2_X1 U293 ( .A1(n116), .A2(n139), .ZN(ab_3__3_) );
  NOR2_X1 U294 ( .A1(n117), .A2(n139), .ZN(ab_3__2_) );
  NOR2_X1 U295 ( .A1(n99), .A2(n139), .ZN(ab_3__22_) );
  NOR2_X1 U296 ( .A1(n96), .A2(n139), .ZN(ab_3__21_) );
  NOR2_X1 U297 ( .A1(n100), .A2(n139), .ZN(ab_3__20_) );
  NOR2_X1 U298 ( .A1(n118), .A2(n139), .ZN(ab_3__1_) );
  NOR2_X1 U299 ( .A1(n90), .A2(n139), .ZN(ab_3__19_) );
  NOR2_X1 U300 ( .A1(n94), .A2(n139), .ZN(ab_3__18_) );
  NOR2_X1 U301 ( .A1(n92), .A2(n139), .ZN(ab_3__17_) );
  NOR2_X1 U302 ( .A1(n103), .A2(n139), .ZN(ab_3__16_) );
  NOR2_X1 U303 ( .A1(n104), .A2(n139), .ZN(ab_3__15_) );
  NOR2_X1 U304 ( .A1(n105), .A2(n139), .ZN(ab_3__14_) );
  NOR2_X1 U305 ( .A1(n106), .A2(n139), .ZN(ab_3__13_) );
  NOR2_X1 U306 ( .A1(n107), .A2(n139), .ZN(ab_3__12_) );
  NOR2_X1 U307 ( .A1(n108), .A2(n139), .ZN(ab_3__11_) );
  NOR2_X1 U308 ( .A1(n109), .A2(n139), .ZN(ab_3__10_) );
  NOR2_X1 U309 ( .A1(n119), .A2(n139), .ZN(ab_3__0_) );
  NOR2_X1 U310 ( .A1(n110), .A2(n140), .ZN(ab_2__9_) );
  NOR2_X1 U311 ( .A1(n111), .A2(n140), .ZN(ab_2__8_) );
  NOR2_X1 U312 ( .A1(n112), .A2(n140), .ZN(ab_2__7_) );
  NOR2_X1 U313 ( .A1(n113), .A2(n140), .ZN(ab_2__6_) );
  NOR2_X1 U314 ( .A1(n114), .A2(n140), .ZN(ab_2__5_) );
  NOR2_X1 U315 ( .A1(n115), .A2(n140), .ZN(ab_2__4_) );
  NOR2_X1 U316 ( .A1(n116), .A2(n140), .ZN(ab_2__3_) );
  NOR2_X1 U317 ( .A1(n117), .A2(n140), .ZN(ab_2__2_) );
  NOR2_X1 U318 ( .A1(n99), .A2(n140), .ZN(ab_2__22_) );
  NOR2_X1 U319 ( .A1(n96), .A2(n140), .ZN(ab_2__21_) );
  NOR2_X1 U320 ( .A1(n100), .A2(n140), .ZN(ab_2__20_) );
  NOR2_X1 U321 ( .A1(n118), .A2(n140), .ZN(ab_2__1_) );
  NOR2_X1 U322 ( .A1(n90), .A2(n140), .ZN(ab_2__19_) );
  NOR2_X1 U323 ( .A1(n94), .A2(n140), .ZN(ab_2__18_) );
  NOR2_X1 U324 ( .A1(n92), .A2(n140), .ZN(ab_2__17_) );
  NOR2_X1 U325 ( .A1(n103), .A2(n140), .ZN(ab_2__16_) );
  NOR2_X1 U326 ( .A1(n104), .A2(n140), .ZN(ab_2__15_) );
  NOR2_X1 U327 ( .A1(n105), .A2(n140), .ZN(ab_2__14_) );
  NOR2_X1 U328 ( .A1(n106), .A2(n140), .ZN(ab_2__13_) );
  NOR2_X1 U329 ( .A1(n107), .A2(n140), .ZN(ab_2__12_) );
  NOR2_X1 U330 ( .A1(n108), .A2(n140), .ZN(ab_2__11_) );
  NOR2_X1 U331 ( .A1(n109), .A2(n140), .ZN(ab_2__10_) );
  NOR2_X1 U332 ( .A1(n119), .A2(n140), .ZN(ab_2__0_) );
  NOR2_X1 U333 ( .A1(n110), .A2(n120), .ZN(ab_22__9_) );
  NOR2_X1 U334 ( .A1(n111), .A2(n120), .ZN(ab_22__8_) );
  NOR2_X1 U335 ( .A1(n112), .A2(n120), .ZN(ab_22__7_) );
  NOR2_X1 U336 ( .A1(n113), .A2(n120), .ZN(ab_22__6_) );
  NOR2_X1 U337 ( .A1(n114), .A2(n120), .ZN(ab_22__5_) );
  NOR2_X1 U338 ( .A1(n115), .A2(n120), .ZN(ab_22__4_) );
  NOR2_X1 U339 ( .A1(n116), .A2(n120), .ZN(ab_22__3_) );
  NOR2_X1 U340 ( .A1(n117), .A2(n120), .ZN(ab_22__2_) );
  NOR2_X1 U341 ( .A1(n99), .A2(n120), .ZN(ab_22__22_) );
  NOR2_X1 U342 ( .A1(n96), .A2(n120), .ZN(ab_22__21_) );
  NOR2_X1 U343 ( .A1(n100), .A2(n120), .ZN(ab_22__20_) );
  NOR2_X1 U344 ( .A1(n118), .A2(n120), .ZN(ab_22__1_) );
  NOR2_X1 U345 ( .A1(n90), .A2(n120), .ZN(ab_22__19_) );
  NOR2_X1 U346 ( .A1(n94), .A2(n120), .ZN(ab_22__18_) );
  NOR2_X1 U347 ( .A1(n92), .A2(n120), .ZN(ab_22__17_) );
  NOR2_X1 U348 ( .A1(n103), .A2(n120), .ZN(ab_22__16_) );
  NOR2_X1 U349 ( .A1(n104), .A2(n120), .ZN(ab_22__15_) );
  NOR2_X1 U350 ( .A1(n105), .A2(n120), .ZN(ab_22__14_) );
  NOR2_X1 U351 ( .A1(n106), .A2(n120), .ZN(ab_22__13_) );
  NOR2_X1 U352 ( .A1(n107), .A2(n120), .ZN(ab_22__12_) );
  NOR2_X1 U353 ( .A1(n108), .A2(n120), .ZN(ab_22__11_) );
  NOR2_X1 U354 ( .A1(n109), .A2(n120), .ZN(ab_22__10_) );
  NOR2_X1 U355 ( .A1(n119), .A2(n120), .ZN(ab_22__0_) );
  NOR2_X1 U356 ( .A1(n110), .A2(n121), .ZN(ab_21__9_) );
  NOR2_X1 U357 ( .A1(n111), .A2(n121), .ZN(ab_21__8_) );
  NOR2_X1 U358 ( .A1(n112), .A2(n121), .ZN(ab_21__7_) );
  NOR2_X1 U359 ( .A1(n113), .A2(n121), .ZN(ab_21__6_) );
  NOR2_X1 U360 ( .A1(n114), .A2(n121), .ZN(ab_21__5_) );
  NOR2_X1 U361 ( .A1(n115), .A2(n121), .ZN(ab_21__4_) );
  NOR2_X1 U362 ( .A1(n116), .A2(n121), .ZN(ab_21__3_) );
  NOR2_X1 U363 ( .A1(n117), .A2(n121), .ZN(ab_21__2_) );
  NOR2_X1 U364 ( .A1(n99), .A2(n121), .ZN(ab_21__22_) );
  NOR2_X1 U365 ( .A1(n96), .A2(n121), .ZN(ab_21__21_) );
  NOR2_X1 U366 ( .A1(n100), .A2(n121), .ZN(ab_21__20_) );
  NOR2_X1 U367 ( .A1(n118), .A2(n121), .ZN(ab_21__1_) );
  NOR2_X1 U368 ( .A1(n90), .A2(n121), .ZN(ab_21__19_) );
  NOR2_X1 U369 ( .A1(n94), .A2(n121), .ZN(ab_21__18_) );
  NOR2_X1 U370 ( .A1(n92), .A2(n121), .ZN(ab_21__17_) );
  NOR2_X1 U371 ( .A1(n103), .A2(n121), .ZN(ab_21__16_) );
  NOR2_X1 U372 ( .A1(n104), .A2(n121), .ZN(ab_21__15_) );
  NOR2_X1 U373 ( .A1(n105), .A2(n121), .ZN(ab_21__14_) );
  NOR2_X1 U374 ( .A1(n106), .A2(n121), .ZN(ab_21__13_) );
  NOR2_X1 U375 ( .A1(n107), .A2(n121), .ZN(ab_21__12_) );
  NOR2_X1 U376 ( .A1(n108), .A2(n121), .ZN(ab_21__11_) );
  NOR2_X1 U377 ( .A1(n109), .A2(n121), .ZN(ab_21__10_) );
  NOR2_X1 U378 ( .A1(n119), .A2(n121), .ZN(ab_21__0_) );
  NOR2_X1 U379 ( .A1(n110), .A2(n122), .ZN(ab_20__9_) );
  NOR2_X1 U380 ( .A1(n111), .A2(n122), .ZN(ab_20__8_) );
  NOR2_X1 U381 ( .A1(n112), .A2(n122), .ZN(ab_20__7_) );
  NOR2_X1 U382 ( .A1(n113), .A2(n122), .ZN(ab_20__6_) );
  NOR2_X1 U383 ( .A1(n114), .A2(n122), .ZN(ab_20__5_) );
  NOR2_X1 U384 ( .A1(n115), .A2(n122), .ZN(ab_20__4_) );
  NOR2_X1 U385 ( .A1(n116), .A2(n122), .ZN(ab_20__3_) );
  NOR2_X1 U386 ( .A1(n117), .A2(n122), .ZN(ab_20__2_) );
  NOR2_X1 U387 ( .A1(n99), .A2(n122), .ZN(ab_20__22_) );
  NOR2_X1 U388 ( .A1(n96), .A2(n122), .ZN(ab_20__21_) );
  NOR2_X1 U389 ( .A1(n100), .A2(n122), .ZN(ab_20__20_) );
  NOR2_X1 U390 ( .A1(n118), .A2(n122), .ZN(ab_20__1_) );
  NOR2_X1 U391 ( .A1(n90), .A2(n122), .ZN(ab_20__19_) );
  NOR2_X1 U392 ( .A1(n94), .A2(n122), .ZN(ab_20__18_) );
  NOR2_X1 U393 ( .A1(n92), .A2(n122), .ZN(ab_20__17_) );
  NOR2_X1 U394 ( .A1(n103), .A2(n122), .ZN(ab_20__16_) );
  NOR2_X1 U395 ( .A1(n104), .A2(n122), .ZN(ab_20__15_) );
  NOR2_X1 U396 ( .A1(n105), .A2(n122), .ZN(ab_20__14_) );
  NOR2_X1 U397 ( .A1(n106), .A2(n122), .ZN(ab_20__13_) );
  NOR2_X1 U398 ( .A1(n107), .A2(n122), .ZN(ab_20__12_) );
  NOR2_X1 U399 ( .A1(n108), .A2(n122), .ZN(ab_20__11_) );
  NOR2_X1 U400 ( .A1(n109), .A2(n122), .ZN(ab_20__10_) );
  NOR2_X1 U401 ( .A1(n119), .A2(n122), .ZN(ab_20__0_) );
  NOR2_X1 U402 ( .A1(n110), .A2(n97), .ZN(ab_1__9_) );
  NOR2_X1 U403 ( .A1(n111), .A2(n97), .ZN(ab_1__8_) );
  NOR2_X1 U404 ( .A1(n112), .A2(n97), .ZN(ab_1__7_) );
  NOR2_X1 U405 ( .A1(n113), .A2(n97), .ZN(ab_1__6_) );
  NOR2_X1 U406 ( .A1(n114), .A2(n97), .ZN(ab_1__5_) );
  NOR2_X1 U407 ( .A1(n115), .A2(n97), .ZN(ab_1__4_) );
  NOR2_X1 U408 ( .A1(n116), .A2(n97), .ZN(ab_1__3_) );
  NOR2_X1 U409 ( .A1(n117), .A2(n97), .ZN(ab_1__2_) );
  NOR2_X1 U410 ( .A1(n99), .A2(n97), .ZN(ab_1__22_) );
  NOR2_X1 U411 ( .A1(n94), .A2(n97), .ZN(ab_1__18_) );
  NOR2_X1 U412 ( .A1(n91), .A2(n97), .ZN(ab_1__17_) );
  NOR2_X1 U413 ( .A1(n103), .A2(n97), .ZN(ab_1__16_) );
  NOR2_X1 U414 ( .A1(n104), .A2(n97), .ZN(ab_1__15_) );
  NOR2_X1 U415 ( .A1(n105), .A2(n97), .ZN(ab_1__14_) );
  NOR2_X1 U416 ( .A1(n106), .A2(n97), .ZN(ab_1__13_) );
  NOR2_X1 U417 ( .A1(n107), .A2(n97), .ZN(ab_1__12_) );
  NOR2_X1 U418 ( .A1(n108), .A2(n97), .ZN(ab_1__11_) );
  NOR2_X1 U419 ( .A1(n109), .A2(n97), .ZN(ab_1__10_) );
  NOR2_X1 U420 ( .A1(n110), .A2(n123), .ZN(ab_19__9_) );
  NOR2_X1 U421 ( .A1(n111), .A2(n123), .ZN(ab_19__8_) );
  NOR2_X1 U422 ( .A1(n112), .A2(n123), .ZN(ab_19__7_) );
  NOR2_X1 U423 ( .A1(n113), .A2(n123), .ZN(ab_19__6_) );
  NOR2_X1 U424 ( .A1(n114), .A2(n123), .ZN(ab_19__5_) );
  NOR2_X1 U425 ( .A1(n115), .A2(n123), .ZN(ab_19__4_) );
  NOR2_X1 U426 ( .A1(n116), .A2(n123), .ZN(ab_19__3_) );
  NOR2_X1 U427 ( .A1(n117), .A2(n123), .ZN(ab_19__2_) );
  NOR2_X1 U428 ( .A1(n99), .A2(n123), .ZN(ab_19__22_) );
  NOR2_X1 U429 ( .A1(n96), .A2(n123), .ZN(ab_19__21_) );
  NOR2_X1 U430 ( .A1(n100), .A2(n123), .ZN(ab_19__20_) );
  NOR2_X1 U431 ( .A1(n118), .A2(n123), .ZN(ab_19__1_) );
  NOR2_X1 U432 ( .A1(n90), .A2(n123), .ZN(ab_19__19_) );
  NOR2_X1 U433 ( .A1(n94), .A2(n123), .ZN(ab_19__18_) );
  NOR2_X1 U434 ( .A1(n92), .A2(n123), .ZN(ab_19__17_) );
  NOR2_X1 U435 ( .A1(n103), .A2(n123), .ZN(ab_19__16_) );
  NOR2_X1 U436 ( .A1(n104), .A2(n123), .ZN(ab_19__15_) );
  NOR2_X1 U437 ( .A1(n105), .A2(n123), .ZN(ab_19__14_) );
  NOR2_X1 U438 ( .A1(n106), .A2(n123), .ZN(ab_19__13_) );
  NOR2_X1 U439 ( .A1(n107), .A2(n123), .ZN(ab_19__12_) );
  NOR2_X1 U440 ( .A1(n108), .A2(n123), .ZN(ab_19__11_) );
  NOR2_X1 U441 ( .A1(n109), .A2(n123), .ZN(ab_19__10_) );
  NOR2_X1 U442 ( .A1(n119), .A2(n123), .ZN(ab_19__0_) );
  NOR2_X1 U443 ( .A1(n110), .A2(n124), .ZN(ab_18__9_) );
  NOR2_X1 U444 ( .A1(n111), .A2(n124), .ZN(ab_18__8_) );
  NOR2_X1 U445 ( .A1(n112), .A2(n124), .ZN(ab_18__7_) );
  NOR2_X1 U446 ( .A1(n113), .A2(n124), .ZN(ab_18__6_) );
  NOR2_X1 U447 ( .A1(n114), .A2(n124), .ZN(ab_18__5_) );
  NOR2_X1 U448 ( .A1(n115), .A2(n124), .ZN(ab_18__4_) );
  NOR2_X1 U449 ( .A1(n116), .A2(n124), .ZN(ab_18__3_) );
  NOR2_X1 U450 ( .A1(n117), .A2(n124), .ZN(ab_18__2_) );
  NOR2_X1 U451 ( .A1(n99), .A2(n124), .ZN(ab_18__22_) );
  NOR2_X1 U452 ( .A1(n96), .A2(n124), .ZN(ab_18__21_) );
  NOR2_X1 U453 ( .A1(n100), .A2(n124), .ZN(ab_18__20_) );
  NOR2_X1 U454 ( .A1(n118), .A2(n124), .ZN(ab_18__1_) );
  NOR2_X1 U455 ( .A1(n90), .A2(n124), .ZN(ab_18__19_) );
  NOR2_X1 U456 ( .A1(n94), .A2(n124), .ZN(ab_18__18_) );
  NOR2_X1 U457 ( .A1(n92), .A2(n124), .ZN(ab_18__17_) );
  NOR2_X1 U458 ( .A1(n103), .A2(n124), .ZN(ab_18__16_) );
  NOR2_X1 U459 ( .A1(n104), .A2(n124), .ZN(ab_18__15_) );
  NOR2_X1 U460 ( .A1(n105), .A2(n124), .ZN(ab_18__14_) );
  NOR2_X1 U461 ( .A1(n106), .A2(n124), .ZN(ab_18__13_) );
  NOR2_X1 U462 ( .A1(n107), .A2(n124), .ZN(ab_18__12_) );
  NOR2_X1 U463 ( .A1(n108), .A2(n124), .ZN(ab_18__11_) );
  NOR2_X1 U464 ( .A1(n109), .A2(n124), .ZN(ab_18__10_) );
  NOR2_X1 U465 ( .A1(n119), .A2(n124), .ZN(ab_18__0_) );
  NOR2_X1 U466 ( .A1(n110), .A2(n125), .ZN(ab_17__9_) );
  NOR2_X1 U467 ( .A1(n111), .A2(n125), .ZN(ab_17__8_) );
  NOR2_X1 U468 ( .A1(n112), .A2(n125), .ZN(ab_17__7_) );
  NOR2_X1 U469 ( .A1(n113), .A2(n125), .ZN(ab_17__6_) );
  NOR2_X1 U470 ( .A1(n114), .A2(n125), .ZN(ab_17__5_) );
  NOR2_X1 U471 ( .A1(n115), .A2(n125), .ZN(ab_17__4_) );
  NOR2_X1 U472 ( .A1(n116), .A2(n125), .ZN(ab_17__3_) );
  NOR2_X1 U473 ( .A1(n117), .A2(n125), .ZN(ab_17__2_) );
  NOR2_X1 U474 ( .A1(n99), .A2(n125), .ZN(ab_17__22_) );
  NOR2_X1 U475 ( .A1(n96), .A2(n125), .ZN(ab_17__21_) );
  NOR2_X1 U476 ( .A1(n100), .A2(n125), .ZN(ab_17__20_) );
  NOR2_X1 U477 ( .A1(n118), .A2(n125), .ZN(ab_17__1_) );
  NOR2_X1 U478 ( .A1(n90), .A2(n125), .ZN(ab_17__19_) );
  NOR2_X1 U479 ( .A1(n94), .A2(n125), .ZN(ab_17__18_) );
  NOR2_X1 U480 ( .A1(n92), .A2(n125), .ZN(ab_17__17_) );
  NOR2_X1 U481 ( .A1(n103), .A2(n125), .ZN(ab_17__16_) );
  NOR2_X1 U482 ( .A1(n104), .A2(n125), .ZN(ab_17__15_) );
  NOR2_X1 U483 ( .A1(n105), .A2(n125), .ZN(ab_17__14_) );
  NOR2_X1 U484 ( .A1(n106), .A2(n125), .ZN(ab_17__13_) );
  NOR2_X1 U485 ( .A1(n107), .A2(n125), .ZN(ab_17__12_) );
  NOR2_X1 U486 ( .A1(n108), .A2(n125), .ZN(ab_17__11_) );
  NOR2_X1 U487 ( .A1(n109), .A2(n125), .ZN(ab_17__10_) );
  NOR2_X1 U488 ( .A1(n119), .A2(n125), .ZN(ab_17__0_) );
  NOR2_X1 U489 ( .A1(n110), .A2(n126), .ZN(ab_16__9_) );
  NOR2_X1 U490 ( .A1(n111), .A2(n126), .ZN(ab_16__8_) );
  NOR2_X1 U491 ( .A1(n112), .A2(n126), .ZN(ab_16__7_) );
  NOR2_X1 U492 ( .A1(n113), .A2(n126), .ZN(ab_16__6_) );
  NOR2_X1 U493 ( .A1(n114), .A2(n126), .ZN(ab_16__5_) );
  NOR2_X1 U494 ( .A1(n115), .A2(n126), .ZN(ab_16__4_) );
  NOR2_X1 U495 ( .A1(n116), .A2(n126), .ZN(ab_16__3_) );
  NOR2_X1 U496 ( .A1(n117), .A2(n126), .ZN(ab_16__2_) );
  NOR2_X1 U497 ( .A1(n99), .A2(n126), .ZN(ab_16__22_) );
  NOR2_X1 U498 ( .A1(n96), .A2(n126), .ZN(ab_16__21_) );
  NOR2_X1 U499 ( .A1(n100), .A2(n126), .ZN(ab_16__20_) );
  NOR2_X1 U500 ( .A1(n118), .A2(n126), .ZN(ab_16__1_) );
  NOR2_X1 U501 ( .A1(n90), .A2(n126), .ZN(ab_16__19_) );
  NOR2_X1 U502 ( .A1(n94), .A2(n126), .ZN(ab_16__18_) );
  NOR2_X1 U503 ( .A1(n92), .A2(n126), .ZN(ab_16__17_) );
  NOR2_X1 U504 ( .A1(n103), .A2(n126), .ZN(ab_16__16_) );
  NOR2_X1 U505 ( .A1(n104), .A2(n126), .ZN(ab_16__15_) );
  NOR2_X1 U506 ( .A1(n105), .A2(n126), .ZN(ab_16__14_) );
  NOR2_X1 U507 ( .A1(n106), .A2(n126), .ZN(ab_16__13_) );
  NOR2_X1 U508 ( .A1(n107), .A2(n126), .ZN(ab_16__12_) );
  NOR2_X1 U509 ( .A1(n108), .A2(n126), .ZN(ab_16__11_) );
  NOR2_X1 U510 ( .A1(n109), .A2(n126), .ZN(ab_16__10_) );
  NOR2_X1 U511 ( .A1(n119), .A2(n126), .ZN(ab_16__0_) );
  NOR2_X1 U512 ( .A1(n110), .A2(n127), .ZN(ab_15__9_) );
  NOR2_X1 U513 ( .A1(n111), .A2(n127), .ZN(ab_15__8_) );
  NOR2_X1 U514 ( .A1(n112), .A2(n127), .ZN(ab_15__7_) );
  NOR2_X1 U515 ( .A1(n113), .A2(n127), .ZN(ab_15__6_) );
  NOR2_X1 U516 ( .A1(n114), .A2(n127), .ZN(ab_15__5_) );
  NOR2_X1 U517 ( .A1(n115), .A2(n127), .ZN(ab_15__4_) );
  NOR2_X1 U518 ( .A1(n116), .A2(n127), .ZN(ab_15__3_) );
  NOR2_X1 U519 ( .A1(n117), .A2(n127), .ZN(ab_15__2_) );
  NOR2_X1 U520 ( .A1(n99), .A2(n127), .ZN(ab_15__22_) );
  NOR2_X1 U521 ( .A1(n96), .A2(n127), .ZN(ab_15__21_) );
  NOR2_X1 U522 ( .A1(n100), .A2(n127), .ZN(ab_15__20_) );
  NOR2_X1 U523 ( .A1(n118), .A2(n127), .ZN(ab_15__1_) );
  NOR2_X1 U524 ( .A1(n90), .A2(n127), .ZN(ab_15__19_) );
  NOR2_X1 U525 ( .A1(n94), .A2(n127), .ZN(ab_15__18_) );
  NOR2_X1 U526 ( .A1(n92), .A2(n127), .ZN(ab_15__17_) );
  NOR2_X1 U527 ( .A1(n103), .A2(n127), .ZN(ab_15__16_) );
  NOR2_X1 U528 ( .A1(n104), .A2(n127), .ZN(ab_15__15_) );
  NOR2_X1 U529 ( .A1(n105), .A2(n127), .ZN(ab_15__14_) );
  NOR2_X1 U530 ( .A1(n106), .A2(n127), .ZN(ab_15__13_) );
  NOR2_X1 U531 ( .A1(n107), .A2(n127), .ZN(ab_15__12_) );
  NOR2_X1 U532 ( .A1(n108), .A2(n127), .ZN(ab_15__11_) );
  NOR2_X1 U533 ( .A1(n109), .A2(n127), .ZN(ab_15__10_) );
  NOR2_X1 U534 ( .A1(n119), .A2(n127), .ZN(ab_15__0_) );
  NOR2_X1 U535 ( .A1(n110), .A2(n128), .ZN(ab_14__9_) );
  NOR2_X1 U536 ( .A1(n111), .A2(n128), .ZN(ab_14__8_) );
  NOR2_X1 U537 ( .A1(n112), .A2(n128), .ZN(ab_14__7_) );
  NOR2_X1 U538 ( .A1(n113), .A2(n128), .ZN(ab_14__6_) );
  NOR2_X1 U539 ( .A1(n114), .A2(n128), .ZN(ab_14__5_) );
  NOR2_X1 U540 ( .A1(n115), .A2(n128), .ZN(ab_14__4_) );
  NOR2_X1 U541 ( .A1(n116), .A2(n128), .ZN(ab_14__3_) );
  NOR2_X1 U542 ( .A1(n117), .A2(n128), .ZN(ab_14__2_) );
  NOR2_X1 U543 ( .A1(n99), .A2(n128), .ZN(ab_14__22_) );
  NOR2_X1 U544 ( .A1(n96), .A2(n128), .ZN(ab_14__21_) );
  NOR2_X1 U545 ( .A1(n100), .A2(n128), .ZN(ab_14__20_) );
  NOR2_X1 U546 ( .A1(n118), .A2(n128), .ZN(ab_14__1_) );
  NOR2_X1 U547 ( .A1(n90), .A2(n128), .ZN(ab_14__19_) );
  NOR2_X1 U548 ( .A1(n94), .A2(n128), .ZN(ab_14__18_) );
  NOR2_X1 U549 ( .A1(n92), .A2(n128), .ZN(ab_14__17_) );
  NOR2_X1 U550 ( .A1(n103), .A2(n128), .ZN(ab_14__16_) );
  NOR2_X1 U551 ( .A1(n104), .A2(n128), .ZN(ab_14__15_) );
  NOR2_X1 U552 ( .A1(n105), .A2(n128), .ZN(ab_14__14_) );
  NOR2_X1 U553 ( .A1(n106), .A2(n128), .ZN(ab_14__13_) );
  NOR2_X1 U554 ( .A1(n107), .A2(n128), .ZN(ab_14__12_) );
  NOR2_X1 U555 ( .A1(n108), .A2(n128), .ZN(ab_14__11_) );
  NOR2_X1 U556 ( .A1(n109), .A2(n128), .ZN(ab_14__10_) );
  NOR2_X1 U557 ( .A1(n119), .A2(n128), .ZN(ab_14__0_) );
  NOR2_X1 U558 ( .A1(n110), .A2(n129), .ZN(ab_13__9_) );
  NOR2_X1 U559 ( .A1(n111), .A2(n129), .ZN(ab_13__8_) );
  NOR2_X1 U560 ( .A1(n112), .A2(n129), .ZN(ab_13__7_) );
  NOR2_X1 U561 ( .A1(n113), .A2(n129), .ZN(ab_13__6_) );
  NOR2_X1 U562 ( .A1(n114), .A2(n129), .ZN(ab_13__5_) );
  NOR2_X1 U563 ( .A1(n115), .A2(n129), .ZN(ab_13__4_) );
  NOR2_X1 U564 ( .A1(n116), .A2(n129), .ZN(ab_13__3_) );
  NOR2_X1 U565 ( .A1(n117), .A2(n129), .ZN(ab_13__2_) );
  NOR2_X1 U566 ( .A1(n99), .A2(n129), .ZN(ab_13__22_) );
  NOR2_X1 U567 ( .A1(n96), .A2(n129), .ZN(ab_13__21_) );
  NOR2_X1 U568 ( .A1(n100), .A2(n129), .ZN(ab_13__20_) );
  NOR2_X1 U569 ( .A1(n118), .A2(n129), .ZN(ab_13__1_) );
  NOR2_X1 U570 ( .A1(n90), .A2(n129), .ZN(ab_13__19_) );
  NOR2_X1 U571 ( .A1(n94), .A2(n129), .ZN(ab_13__18_) );
  NOR2_X1 U572 ( .A1(n92), .A2(n129), .ZN(ab_13__17_) );
  NOR2_X1 U573 ( .A1(n103), .A2(n129), .ZN(ab_13__16_) );
  NOR2_X1 U574 ( .A1(n104), .A2(n129), .ZN(ab_13__15_) );
  NOR2_X1 U575 ( .A1(n105), .A2(n129), .ZN(ab_13__14_) );
  NOR2_X1 U576 ( .A1(n106), .A2(n129), .ZN(ab_13__13_) );
  NOR2_X1 U577 ( .A1(n107), .A2(n129), .ZN(ab_13__12_) );
  NOR2_X1 U578 ( .A1(n108), .A2(n129), .ZN(ab_13__11_) );
  NOR2_X1 U579 ( .A1(n109), .A2(n129), .ZN(ab_13__10_) );
  NOR2_X1 U580 ( .A1(n119), .A2(n129), .ZN(ab_13__0_) );
  NOR2_X1 U581 ( .A1(n110), .A2(n130), .ZN(ab_12__9_) );
  NOR2_X1 U582 ( .A1(n111), .A2(n130), .ZN(ab_12__8_) );
  NOR2_X1 U583 ( .A1(n112), .A2(n130), .ZN(ab_12__7_) );
  NOR2_X1 U584 ( .A1(n113), .A2(n130), .ZN(ab_12__6_) );
  NOR2_X1 U585 ( .A1(n114), .A2(n130), .ZN(ab_12__5_) );
  NOR2_X1 U586 ( .A1(n115), .A2(n130), .ZN(ab_12__4_) );
  NOR2_X1 U587 ( .A1(n116), .A2(n130), .ZN(ab_12__3_) );
  NOR2_X1 U588 ( .A1(n117), .A2(n130), .ZN(ab_12__2_) );
  NOR2_X1 U589 ( .A1(n99), .A2(n130), .ZN(ab_12__22_) );
  NOR2_X1 U590 ( .A1(n96), .A2(n130), .ZN(ab_12__21_) );
  NOR2_X1 U591 ( .A1(n100), .A2(n130), .ZN(ab_12__20_) );
  NOR2_X1 U592 ( .A1(n118), .A2(n130), .ZN(ab_12__1_) );
  NOR2_X1 U593 ( .A1(n90), .A2(n130), .ZN(ab_12__19_) );
  NOR2_X1 U594 ( .A1(n94), .A2(n130), .ZN(ab_12__18_) );
  NOR2_X1 U595 ( .A1(n92), .A2(n130), .ZN(ab_12__17_) );
  NOR2_X1 U596 ( .A1(n103), .A2(n130), .ZN(ab_12__16_) );
  NOR2_X1 U597 ( .A1(n104), .A2(n130), .ZN(ab_12__15_) );
  NOR2_X1 U598 ( .A1(n105), .A2(n130), .ZN(ab_12__14_) );
  NOR2_X1 U599 ( .A1(n106), .A2(n130), .ZN(ab_12__13_) );
  NOR2_X1 U600 ( .A1(n107), .A2(n130), .ZN(ab_12__12_) );
  NOR2_X1 U601 ( .A1(n108), .A2(n130), .ZN(ab_12__11_) );
  NOR2_X1 U602 ( .A1(n109), .A2(n130), .ZN(ab_12__10_) );
  NOR2_X1 U603 ( .A1(n119), .A2(n130), .ZN(ab_12__0_) );
  NOR2_X1 U604 ( .A1(n110), .A2(n131), .ZN(ab_11__9_) );
  NOR2_X1 U605 ( .A1(n111), .A2(n131), .ZN(ab_11__8_) );
  NOR2_X1 U606 ( .A1(n112), .A2(n131), .ZN(ab_11__7_) );
  NOR2_X1 U607 ( .A1(n113), .A2(n131), .ZN(ab_11__6_) );
  NOR2_X1 U608 ( .A1(n114), .A2(n131), .ZN(ab_11__5_) );
  NOR2_X1 U609 ( .A1(n115), .A2(n131), .ZN(ab_11__4_) );
  NOR2_X1 U610 ( .A1(n116), .A2(n131), .ZN(ab_11__3_) );
  NOR2_X1 U611 ( .A1(n117), .A2(n131), .ZN(ab_11__2_) );
  NOR2_X1 U612 ( .A1(n99), .A2(n131), .ZN(ab_11__22_) );
  NOR2_X1 U613 ( .A1(n96), .A2(n131), .ZN(ab_11__21_) );
  NOR2_X1 U614 ( .A1(n100), .A2(n131), .ZN(ab_11__20_) );
  NOR2_X1 U615 ( .A1(n118), .A2(n131), .ZN(ab_11__1_) );
  NOR2_X1 U616 ( .A1(n90), .A2(n131), .ZN(ab_11__19_) );
  NOR2_X1 U617 ( .A1(n94), .A2(n131), .ZN(ab_11__18_) );
  NOR2_X1 U618 ( .A1(n92), .A2(n131), .ZN(ab_11__17_) );
  NOR2_X1 U619 ( .A1(n103), .A2(n131), .ZN(ab_11__16_) );
  NOR2_X1 U620 ( .A1(n104), .A2(n131), .ZN(ab_11__15_) );
  NOR2_X1 U621 ( .A1(n105), .A2(n131), .ZN(ab_11__14_) );
  NOR2_X1 U622 ( .A1(n106), .A2(n131), .ZN(ab_11__13_) );
  NOR2_X1 U623 ( .A1(n107), .A2(n131), .ZN(ab_11__12_) );
  NOR2_X1 U624 ( .A1(n108), .A2(n131), .ZN(ab_11__11_) );
  NOR2_X1 U625 ( .A1(n109), .A2(n131), .ZN(ab_11__10_) );
  NOR2_X1 U626 ( .A1(n119), .A2(n131), .ZN(ab_11__0_) );
  NOR2_X1 U627 ( .A1(n110), .A2(n132), .ZN(ab_10__9_) );
  NOR2_X1 U628 ( .A1(n111), .A2(n132), .ZN(ab_10__8_) );
  NOR2_X1 U629 ( .A1(n112), .A2(n132), .ZN(ab_10__7_) );
  NOR2_X1 U630 ( .A1(n113), .A2(n132), .ZN(ab_10__6_) );
  NOR2_X1 U631 ( .A1(n114), .A2(n132), .ZN(ab_10__5_) );
  NOR2_X1 U632 ( .A1(n115), .A2(n132), .ZN(ab_10__4_) );
  NOR2_X1 U633 ( .A1(n116), .A2(n132), .ZN(ab_10__3_) );
  NOR2_X1 U634 ( .A1(n117), .A2(n132), .ZN(ab_10__2_) );
  NOR2_X1 U635 ( .A1(n99), .A2(n132), .ZN(ab_10__22_) );
  NOR2_X1 U636 ( .A1(n96), .A2(n132), .ZN(ab_10__21_) );
  NOR2_X1 U637 ( .A1(n100), .A2(n132), .ZN(ab_10__20_) );
  NOR2_X1 U638 ( .A1(n118), .A2(n132), .ZN(ab_10__1_) );
  NOR2_X1 U639 ( .A1(n90), .A2(n132), .ZN(ab_10__19_) );
  NOR2_X1 U640 ( .A1(n94), .A2(n132), .ZN(ab_10__18_) );
  NOR2_X1 U641 ( .A1(n92), .A2(n132), .ZN(ab_10__17_) );
  NOR2_X1 U642 ( .A1(n103), .A2(n132), .ZN(ab_10__16_) );
  NOR2_X1 U643 ( .A1(n104), .A2(n132), .ZN(ab_10__15_) );
  NOR2_X1 U644 ( .A1(n105), .A2(n132), .ZN(ab_10__14_) );
  NOR2_X1 U645 ( .A1(n106), .A2(n132), .ZN(ab_10__13_) );
  NOR2_X1 U646 ( .A1(n107), .A2(n132), .ZN(ab_10__12_) );
  NOR2_X1 U647 ( .A1(n108), .A2(n132), .ZN(ab_10__11_) );
  NOR2_X1 U648 ( .A1(n109), .A2(n132), .ZN(ab_10__10_) );
  NOR2_X1 U649 ( .A1(n119), .A2(n132), .ZN(ab_10__0_) );
  NOR2_X1 U650 ( .A1(n110), .A2(n141), .ZN(ab_0__9_) );
  NOR2_X1 U651 ( .A1(n111), .A2(n93), .ZN(ab_0__8_) );
  NOR2_X1 U652 ( .A1(n112), .A2(n93), .ZN(ab_0__7_) );
  NOR2_X1 U653 ( .A1(n113), .A2(n93), .ZN(ab_0__6_) );
  NOR2_X1 U654 ( .A1(n114), .A2(n93), .ZN(ab_0__5_) );
  NOR2_X1 U655 ( .A1(n115), .A2(n93), .ZN(ab_0__4_) );
  NOR2_X1 U656 ( .A1(n116), .A2(n93), .ZN(ab_0__3_) );
  NOR2_X1 U657 ( .A1(n117), .A2(n93), .ZN(ab_0__2_) );
  NOR2_X1 U658 ( .A1(n101), .A2(n141), .ZN(ab_0__19_) );
  NOR2_X1 U659 ( .A1(n94), .A2(n141), .ZN(ab_0__18_) );
  NOR2_X1 U660 ( .A1(n91), .A2(n141), .ZN(ab_0__17_) );
  NOR2_X1 U661 ( .A1(n103), .A2(n141), .ZN(ab_0__16_) );
  NOR2_X1 U662 ( .A1(n104), .A2(n141), .ZN(ab_0__15_) );
  NOR2_X1 U663 ( .A1(n105), .A2(n141), .ZN(ab_0__14_) );
  NOR2_X1 U664 ( .A1(n106), .A2(n141), .ZN(ab_0__13_) );
  NOR2_X1 U665 ( .A1(n107), .A2(n141), .ZN(ab_0__12_) );
  NOR2_X1 U666 ( .A1(n108), .A2(n141), .ZN(ab_0__11_) );
  NOR2_X1 U667 ( .A1(n109), .A2(n141), .ZN(ab_0__10_) );
  AND3_X1 U668 ( .A1(ab_1__1_), .A2(B[0]), .A3(n95), .ZN(CARRYB_1__0_) );
  NOR2_X1 U669 ( .A1(n97), .A2(n118), .ZN(ab_1__1_) );
endmodule


module FPM_DW01_add_1 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:2] carry;

  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2_X1 U1 ( .A1(B[0]), .A2(A[0]), .ZN(n1) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module FPM ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [31:0] result;
  wire   N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19,
         N20, N21, N22, N23, N24, N25, N26, N27, N28, N47, N48, N49, N50, N51,
         N52, N53, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n470, n480, n490, n500, n510, n520, n530, n54, n55,
         N31, N30, add_0_root_sub_1_root_add_30_2_A_0_,
         add_0_root_sub_1_root_add_30_2_A_1_,
         add_0_root_sub_1_root_add_30_2_A_2_,
         add_0_root_sub_1_root_add_30_2_A_3_,
         add_0_root_sub_1_root_add_30_2_A_4_,
         add_0_root_sub_1_root_add_30_2_A_5_,
         add_0_root_sub_1_root_add_30_2_A_6_,
         add_0_root_sub_1_root_add_30_2_A_7_, n1, n2, n3, n4, n560, n60, n70,
         n80, n90, n100, n110, n120, n130, n140, n150, n160, n170, n180, n190,
         n200, n210, n220, n230, n240, n250, n260, n270, n280, n29, n300,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16,
         SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18,
         SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20,
         SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22,
         SYNOPSYS_UNCONNECTED_23;
  wire   [7:2] add_0_root_sub_1_root_add_30_2_carry;

  FPM_DW02_mult_0 mult_28 ( .A({1'b1, a[22:0]}), .B({1'b1, b[22:0]}), .TC(1'b0), .PRODUCT({N31, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, 
        N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, 
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, 
        SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, 
        SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, 
        SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23}) );
  FPM_DW01_add_1 add_2_root_sub_1_root_add_30_2 ( .A(b[30:23]), .B(a[30:23]), 
        .CI(1'b0), .SUM({add_0_root_sub_1_root_add_30_2_A_7_, 
        add_0_root_sub_1_root_add_30_2_A_6_, 
        add_0_root_sub_1_root_add_30_2_A_5_, 
        add_0_root_sub_1_root_add_30_2_A_4_, 
        add_0_root_sub_1_root_add_30_2_A_3_, 
        add_0_root_sub_1_root_add_30_2_A_2_, 
        add_0_root_sub_1_root_add_30_2_A_1_, 
        add_0_root_sub_1_root_add_30_2_A_0_}) );
  FA_X1 add_0_root_sub_1_root_add_30_2_U1_1 ( .A(
        add_0_root_sub_1_root_add_30_2_A_1_), .B(n3), .CI(n1), .CO(
        add_0_root_sub_1_root_add_30_2_carry[2]), .S(N47) );
  FA_X1 add_0_root_sub_1_root_add_30_2_U1_6 ( .A(
        add_0_root_sub_1_root_add_30_2_A_6_), .B(1'b0), .CI(
        add_0_root_sub_1_root_add_30_2_carry[6]), .CO(
        add_0_root_sub_1_root_add_30_2_carry[7]), .S(N52) );
  FA_X1 add_0_root_sub_1_root_add_30_2_U1_5 ( .A(
        add_0_root_sub_1_root_add_30_2_A_5_), .B(1'b0), .CI(
        add_0_root_sub_1_root_add_30_2_carry[5]), .CO(
        add_0_root_sub_1_root_add_30_2_carry[6]), .S(N51) );
  FA_X1 add_0_root_sub_1_root_add_30_2_U1_4 ( .A(
        add_0_root_sub_1_root_add_30_2_A_4_), .B(1'b0), .CI(
        add_0_root_sub_1_root_add_30_2_carry[4]), .CO(
        add_0_root_sub_1_root_add_30_2_carry[5]), .S(N50) );
  FA_X1 add_0_root_sub_1_root_add_30_2_U1_3 ( .A(
        add_0_root_sub_1_root_add_30_2_A_3_), .B(1'b0), .CI(
        add_0_root_sub_1_root_add_30_2_carry[3]), .CO(
        add_0_root_sub_1_root_add_30_2_carry[4]), .S(N49) );
  FA_X1 add_0_root_sub_1_root_add_30_2_U1_2 ( .A(
        add_0_root_sub_1_root_add_30_2_A_2_), .B(1'b0), .CI(
        add_0_root_sub_1_root_add_30_2_carry[2]), .CO(
        add_0_root_sub_1_root_add_30_2_carry[3]), .S(N48) );
  INV_X1 U3 ( .A(N6), .ZN(n280) );
  AND2_X1 U4 ( .A1(n2), .A2(n300), .ZN(result[23]) );
  OAI22_X1 U5 ( .A1(n4), .A2(n250), .B1(n560), .B2(n260), .ZN(result[3]) );
  OAI22_X1 U6 ( .A1(n4), .A2(n230), .B1(n560), .B2(n240), .ZN(result[5]) );
  OAI22_X1 U7 ( .A1(n4), .A2(n210), .B1(n560), .B2(n220), .ZN(result[7]) );
  OAI22_X1 U8 ( .A1(n4), .A2(n170), .B1(n560), .B2(n180), .ZN(result[11]) );
  OAI22_X1 U9 ( .A1(n4), .A2(n150), .B1(n560), .B2(n160), .ZN(result[13]) );
  OAI22_X1 U10 ( .A1(n4), .A2(n130), .B1(n560), .B2(n140), .ZN(result[15]) );
  OAI22_X1 U11 ( .A1(n4), .A2(n110), .B1(n560), .B2(n120), .ZN(result[17]) );
  OAI22_X1 U12 ( .A1(n4), .A2(n90), .B1(n560), .B2(n100), .ZN(result[19]) );
  OAI22_X1 U13 ( .A1(n4), .A2(n80), .B1(n560), .B2(n90), .ZN(result[20]) );
  OAI22_X1 U14 ( .A1(n4), .A2(n60), .B1(n560), .B2(n70), .ZN(result[22]) );
  INV_X1 U15 ( .A(N28), .ZN(n60) );
  OAI22_X1 U16 ( .A1(n32), .A2(n260), .B1(n33), .B2(n270), .ZN(result[2]) );
  OAI22_X1 U17 ( .A1(n32), .A2(n240), .B1(n33), .B2(n250), .ZN(result[4]) );
  OAI22_X1 U18 ( .A1(n32), .A2(n220), .B1(n33), .B2(n230), .ZN(result[6]) );
  OAI22_X1 U19 ( .A1(n32), .A2(n190), .B1(n560), .B2(n200), .ZN(result[9]) );
  OAI22_X1 U20 ( .A1(n32), .A2(n180), .B1(n33), .B2(n190), .ZN(result[10]) );
  OAI22_X1 U21 ( .A1(n32), .A2(n160), .B1(n33), .B2(n170), .ZN(result[12]) );
  OAI22_X1 U22 ( .A1(n32), .A2(n140), .B1(n33), .B2(n150), .ZN(result[14]) );
  OAI22_X1 U23 ( .A1(n32), .A2(n120), .B1(n33), .B2(n130), .ZN(result[16]) );
  OAI22_X1 U24 ( .A1(n32), .A2(n100), .B1(n33), .B2(n110), .ZN(result[18]) );
  OAI22_X1 U25 ( .A1(n32), .A2(n70), .B1(n33), .B2(n80), .ZN(result[21]) );
  OAI22_X1 U26 ( .A1(n200), .A2(n4), .B1(n33), .B2(n210), .ZN(result[8]) );
  INV_X1 U27 ( .A(N24), .ZN(n100) );
  INV_X1 U28 ( .A(N26), .ZN(n80) );
  INV_X1 U29 ( .A(N21), .ZN(n130) );
  INV_X1 U30 ( .A(N23), .ZN(n110) );
  INV_X1 U31 ( .A(N25), .ZN(n90) );
  INV_X1 U32 ( .A(N27), .ZN(n70) );
  INV_X1 U33 ( .A(N22), .ZN(n120) );
  INV_X1 U34 ( .A(N20), .ZN(n140) );
  INV_X1 U35 ( .A(N9), .ZN(n250) );
  INV_X1 U36 ( .A(N13), .ZN(n210) );
  INV_X1 U37 ( .A(N15), .ZN(n190) );
  INV_X1 U38 ( .A(N19), .ZN(n150) );
  INV_X1 U39 ( .A(N8), .ZN(n260) );
  INV_X1 U40 ( .A(N10), .ZN(n240) );
  INV_X1 U41 ( .A(N11), .ZN(n230) );
  INV_X1 U42 ( .A(N12), .ZN(n220) );
  INV_X1 U43 ( .A(N16), .ZN(n180) );
  INV_X1 U44 ( .A(N17), .ZN(n170) );
  INV_X1 U45 ( .A(N18), .ZN(n160) );
  INV_X1 U46 ( .A(N14), .ZN(n200) );
  INV_X1 U47 ( .A(N7), .ZN(n270) );
  OAI22_X1 U48 ( .A1(n32), .A2(n270), .B1(n33), .B2(n280), .ZN(result[1]) );
  AND2_X1 U49 ( .A1(N47), .A2(n300), .ZN(result[24]) );
  INV_X1 U50 ( .A(n35), .ZN(n300) );
  OAI22_X1 U51 ( .A1(n4), .A2(n280), .B1(n560), .B2(n29), .ZN(result[0]) );
  INV_X1 U52 ( .A(N5), .ZN(n29) );
  AND2_X1 U53 ( .A1(N30), .A2(add_0_root_sub_1_root_add_30_2_A_0_), .ZN(n1) );
  AND2_X1 U54 ( .A1(N51), .A2(n300), .ZN(result[28]) );
  AND2_X1 U55 ( .A1(N52), .A2(n300), .ZN(result[29]) );
  AND2_X1 U56 ( .A1(N48), .A2(n300), .ZN(result[25]) );
  AND2_X1 U57 ( .A1(N49), .A2(n300), .ZN(result[26]) );
  AND2_X1 U58 ( .A1(N50), .A2(n300), .ZN(result[27]) );
  XOR2_X1 U59 ( .A(N30), .B(add_0_root_sub_1_root_add_30_2_A_0_), .Z(n2) );
  OAI22_X1 U60 ( .A1(n36), .A2(n37), .B1(n38), .B2(n39), .ZN(n35) );
  NAND4_X1 U61 ( .A1(n520), .A2(n530), .A3(n54), .A4(n55), .ZN(n36) );
  NAND4_X1 U62 ( .A1(n44), .A2(n45), .A3(n46), .A4(n470), .ZN(n38) );
  NAND4_X1 U63 ( .A1(n480), .A2(n490), .A3(n500), .A4(n510), .ZN(n37) );
  XNOR2_X1 U64 ( .A(add_0_root_sub_1_root_add_30_2_A_7_), .B(
        add_0_root_sub_1_root_add_30_2_carry[7]), .ZN(N53) );
  NAND4_X1 U65 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n39) );
  NOR4_X1 U66 ( .A1(a[15]), .A2(a[14]), .A3(a[13]), .A4(a[12]), .ZN(n41) );
  NOR4_X1 U67 ( .A1(a[19]), .A2(a[18]), .A3(a[17]), .A4(a[16]), .ZN(n42) );
  NOR4_X1 U68 ( .A1(a[9]), .A2(a[8]), .A3(a[7]), .A4(a[6]), .ZN(n470) );
  NOR4_X1 U69 ( .A1(b[9]), .A2(b[8]), .A3(b[7]), .A4(b[6]), .ZN(n55) );
  NOR4_X1 U70 ( .A1(a[5]), .A2(a[4]), .A3(a[3]), .A4(a[30]), .ZN(n46) );
  NOR4_X1 U71 ( .A1(b[5]), .A2(b[4]), .A3(b[3]), .A4(b[30]), .ZN(n54) );
  NOR4_X1 U72 ( .A1(b[15]), .A2(b[14]), .A3(b[13]), .A4(b[12]), .ZN(n490) );
  NOR4_X1 U73 ( .A1(a[2]), .A2(a[29]), .A3(a[28]), .A4(a[27]), .ZN(n45) );
  NOR4_X1 U74 ( .A1(b[2]), .A2(b[29]), .A3(b[28]), .A4(b[27]), .ZN(n530) );
  NOR4_X1 U75 ( .A1(a[26]), .A2(a[25]), .A3(a[24]), .A4(a[23]), .ZN(n44) );
  NOR4_X1 U76 ( .A1(b[26]), .A2(b[25]), .A3(b[24]), .A4(b[23]), .ZN(n520) );
  NOR3_X1 U77 ( .A1(b[0]), .A2(b[11]), .A3(b[10]), .ZN(n480) );
  NOR2_X1 U78 ( .A1(n34), .A2(n35), .ZN(result[31]) );
  XNOR2_X1 U79 ( .A(b[31]), .B(a[31]), .ZN(n34) );
  CLKBUF_X1 U80 ( .A(N31), .Z(n3) );
  NOR4_X1 U81 ( .A1(b[19]), .A2(b[18]), .A3(b[17]), .A4(b[16]), .ZN(n500) );
  NOR4_X1 U82 ( .A1(a[22]), .A2(a[21]), .A3(a[20]), .A4(a[1]), .ZN(n43) );
  NOR3_X1 U83 ( .A1(a[0]), .A2(a[11]), .A3(a[10]), .ZN(n40) );
  AND2_X1 U84 ( .A1(N53), .A2(n300), .ZN(result[30]) );
  NAND2_X1 U85 ( .A1(n3), .A2(n300), .ZN(n32) );
  OR2_X1 U86 ( .A1(n35), .A2(n3), .ZN(n33) );
  OR2_X1 U87 ( .A1(n35), .A2(n3), .ZN(n560) );
  NAND2_X1 U88 ( .A1(n3), .A2(n300), .ZN(n4) );
  NOR4_X1 U89 ( .A1(b[22]), .A2(b[21]), .A3(b[20]), .A4(b[1]), .ZN(n510) );
  INV_X1 U90 ( .A(N31), .ZN(N30) );
endmodule


module regN_N32_1 ( clk, reset, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, reset;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  DFF_X1 out_reg_31_ ( .D(n32), .CK(clk), .Q(out[31]) );
  DFF_X1 out_reg_23_ ( .D(n31), .CK(clk), .Q(out[23]) );
  DFF_X1 out_reg_21_ ( .D(n30), .CK(clk), .Q(out[21]) );
  DFF_X1 out_reg_18_ ( .D(n29), .CK(clk), .Q(out[18]) );
  DFF_X1 out_reg_16_ ( .D(n28), .CK(clk), .Q(out[16]) );
  DFF_X1 out_reg_14_ ( .D(n27), .CK(clk), .Q(out[14]) );
  DFF_X1 out_reg_12_ ( .D(n26), .CK(clk), .Q(out[12]) );
  DFF_X1 out_reg_10_ ( .D(n25), .CK(clk), .Q(out[10]) );
  DFF_X1 out_reg_6_ ( .D(n24), .CK(clk), .Q(out[6]) );
  DFF_X1 out_reg_4_ ( .D(n23), .CK(clk), .Q(out[4]) );
  DFF_X1 out_reg_2_ ( .D(n22), .CK(clk), .Q(out[2]) );
  DFF_X1 out_reg_1_ ( .D(n21), .CK(clk), .Q(out[1]) );
  DFF_X1 out_reg_9_ ( .D(n20), .CK(clk), .Q(out[9]) );
  DFF_X1 out_reg_22_ ( .D(n19), .CK(clk), .Q(out[22]) );
  DFF_X1 out_reg_20_ ( .D(n18), .CK(clk), .Q(out[20]) );
  DFF_X1 out_reg_19_ ( .D(n17), .CK(clk), .Q(out[19]) );
  DFF_X1 out_reg_17_ ( .D(n16), .CK(clk), .Q(out[17]) );
  DFF_X1 out_reg_15_ ( .D(n15), .CK(clk), .Q(out[15]) );
  DFF_X1 out_reg_13_ ( .D(n14), .CK(clk), .Q(out[13]) );
  DFF_X1 out_reg_11_ ( .D(n13), .CK(clk), .Q(out[11]) );
  DFF_X1 out_reg_7_ ( .D(n12), .CK(clk), .Q(out[7]) );
  DFF_X1 out_reg_5_ ( .D(n11), .CK(clk), .Q(out[5]) );
  DFF_X1 out_reg_3_ ( .D(n10), .CK(clk), .Q(out[3]) );
  DFF_X1 out_reg_0_ ( .D(n9), .CK(clk), .Q(out[0]) );
  DFF_X1 out_reg_8_ ( .D(n8), .CK(clk), .Q(out[8]) );
  DFF_X1 out_reg_24_ ( .D(n7), .CK(clk), .Q(out[24]) );
  DFF_X1 out_reg_25_ ( .D(n6), .CK(clk), .Q(out[25]) );
  DFF_X1 out_reg_26_ ( .D(n5), .CK(clk), .Q(out[26]) );
  DFF_X1 out_reg_27_ ( .D(n4), .CK(clk), .Q(out[27]) );
  DFF_X1 out_reg_28_ ( .D(n3), .CK(clk), .Q(out[28]) );
  DFF_X1 out_reg_29_ ( .D(n2), .CK(clk), .Q(out[29]) );
  DFF_X1 out_reg_30_ ( .D(n1), .CK(clk), .Q(out[30]) );
  AND2_X1 U3 ( .A1(in[30]), .A2(n33), .ZN(n1) );
  AND2_X1 U4 ( .A1(in[29]), .A2(n33), .ZN(n2) );
  AND2_X1 U5 ( .A1(in[28]), .A2(n33), .ZN(n3) );
  AND2_X1 U6 ( .A1(in[27]), .A2(n33), .ZN(n4) );
  AND2_X1 U7 ( .A1(in[26]), .A2(n33), .ZN(n5) );
  AND2_X1 U8 ( .A1(in[25]), .A2(n33), .ZN(n6) );
  AND2_X1 U9 ( .A1(in[24]), .A2(n33), .ZN(n7) );
  AND2_X1 U10 ( .A1(in[8]), .A2(n35), .ZN(n8) );
  AND2_X1 U11 ( .A1(in[0]), .A2(n35), .ZN(n9) );
  AND2_X1 U12 ( .A1(in[3]), .A2(n35), .ZN(n10) );
  AND2_X1 U13 ( .A1(in[5]), .A2(n35), .ZN(n11) );
  AND2_X1 U14 ( .A1(in[7]), .A2(n35), .ZN(n12) );
  AND2_X1 U15 ( .A1(in[11]), .A2(n34), .ZN(n13) );
  AND2_X1 U16 ( .A1(in[13]), .A2(n34), .ZN(n14) );
  AND2_X1 U17 ( .A1(in[15]), .A2(n34), .ZN(n15) );
  AND2_X1 U18 ( .A1(in[17]), .A2(n34), .ZN(n16) );
  AND2_X1 U19 ( .A1(in[19]), .A2(n34), .ZN(n17) );
  AND2_X1 U20 ( .A1(in[20]), .A2(n34), .ZN(n18) );
  AND2_X1 U21 ( .A1(in[22]), .A2(n33), .ZN(n19) );
  AND2_X1 U22 ( .A1(in[9]), .A2(n35), .ZN(n20) );
  AND2_X1 U23 ( .A1(in[1]), .A2(n35), .ZN(n21) );
  AND2_X1 U24 ( .A1(in[2]), .A2(n35), .ZN(n22) );
  AND2_X1 U25 ( .A1(in[4]), .A2(n35), .ZN(n23) );
  AND2_X1 U26 ( .A1(in[6]), .A2(n35), .ZN(n24) );
  AND2_X1 U27 ( .A1(in[10]), .A2(n34), .ZN(n25) );
  AND2_X1 U28 ( .A1(in[12]), .A2(n34), .ZN(n26) );
  AND2_X1 U29 ( .A1(in[14]), .A2(n34), .ZN(n27) );
  AND2_X1 U30 ( .A1(in[16]), .A2(n34), .ZN(n28) );
  AND2_X1 U31 ( .A1(in[18]), .A2(n34), .ZN(n29) );
  AND2_X1 U32 ( .A1(in[21]), .A2(n33), .ZN(n30) );
  AND2_X1 U33 ( .A1(in[23]), .A2(n33), .ZN(n31) );
  AND2_X1 U34 ( .A1(in[31]), .A2(n33), .ZN(n32) );
  BUF_X1 U35 ( .A(n36), .Z(n34) );
  BUF_X1 U36 ( .A(n36), .Z(n33) );
  BUF_X1 U37 ( .A(n36), .Z(n35) );
  INV_X1 U38 ( .A(reset), .ZN(n36) );
endmodule


module FPMSeq ( A, B, clk, reset, result );
  input [31:0] A;
  input [31:0] B;
  output [31:0] result;
  input clk, reset;

  wire   [31:0] AReg;
  wire   [31:0] BReg;
  wire   [31:0] resultReg;

  regN_N32_0 regA ( .clk(clk), .reset(reset), .in(A), .out(AReg) );
  regN_N32_2 regB ( .clk(clk), .reset(reset), .in(B), .out(BReg) );
  FPM multiplier ( .a(AReg), .b(BReg), .result(resultReg) );
  regN_N32_1 outA ( .clk(clk), .reset(reset), .in(resultReg), .out(result) );
endmodule


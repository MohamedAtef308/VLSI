
module regN ( clk, reset, in, out );
  input [31:0] in;
  output [31:0] out;
  input clk, reset;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68;

  DFF_X1 out_reg_9_ ( .D(n65), .CK(clk), .Q(out[9]) );
  DFF_X1 out_reg_8_ ( .D(n64), .CK(clk), .Q(out[8]) );
  DFF_X1 out_reg_7_ ( .D(n63), .CK(clk), .Q(out[7]) );
  DFF_X1 out_reg_6_ ( .D(n62), .CK(clk), .Q(out[6]) );
  DFF_X1 out_reg_5_ ( .D(n61), .CK(clk), .Q(out[5]) );
  DFF_X1 out_reg_4_ ( .D(n60), .CK(clk), .Q(out[4]) );
  DFF_X1 out_reg_3_ ( .D(n59), .CK(clk), .Q(out[3]) );
  DFF_X1 out_reg_2_ ( .D(n58), .CK(clk), .Q(out[2]) );
  DFF_X1 out_reg_1_ ( .D(n57), .CK(clk), .Q(out[1]) );
  DFF_X1 out_reg_0_ ( .D(n56), .CK(clk), .Q(out[0]) );
  DFF_X1 out_reg_31_ ( .D(n55), .CK(clk), .Q(out[31]) );
  DFF_X1 out_reg_30_ ( .D(n54), .CK(clk), .Q(out[30]) );
  DFF_X1 out_reg_29_ ( .D(n53), .CK(clk), .Q(out[29]) );
  DFF_X1 out_reg_28_ ( .D(n52), .CK(clk), .Q(out[28]) );
  DFF_X1 out_reg_27_ ( .D(n51), .CK(clk), .Q(out[27]) );
  DFF_X1 out_reg_26_ ( .D(n50), .CK(clk), .Q(out[26]) );
  DFF_X1 out_reg_25_ ( .D(n49), .CK(clk), .Q(out[25]) );
  DFF_X1 out_reg_24_ ( .D(n48), .CK(clk), .Q(out[24]) );
  DFF_X1 out_reg_23_ ( .D(n47), .CK(clk), .Q(out[23]) );
  DFF_X1 out_reg_22_ ( .D(n46), .CK(clk), .Q(out[22]) );
  DFF_X1 out_reg_21_ ( .D(n45), .CK(clk), .Q(out[21]) );
  DFF_X1 out_reg_20_ ( .D(n44), .CK(clk), .Q(out[20]) );
  DFF_X1 out_reg_19_ ( .D(n43), .CK(clk), .Q(out[19]) );
  DFF_X1 out_reg_18_ ( .D(n42), .CK(clk), .Q(out[18]) );
  DFF_X1 out_reg_17_ ( .D(n41), .CK(clk), .Q(out[17]) );
  DFF_X1 out_reg_16_ ( .D(n40), .CK(clk), .Q(out[16]) );
  DFF_X1 out_reg_15_ ( .D(n39), .CK(clk), .Q(out[15]) );
  DFF_X1 out_reg_14_ ( .D(n38), .CK(clk), .Q(out[14]) );
  DFF_X1 out_reg_13_ ( .D(n37), .CK(clk), .Q(out[13]) );
  DFF_X1 out_reg_12_ ( .D(n36), .CK(clk), .Q(out[12]) );
  DFF_X1 out_reg_11_ ( .D(n35), .CK(clk), .Q(out[11]) );
  DFF_X1 out_reg_10_ ( .D(n34), .CK(clk), .Q(out[10]) );
  AND2_X1 U36 ( .A1(in[10]), .A2(n67), .ZN(n34) );
  AND2_X1 U37 ( .A1(in[11]), .A2(n67), .ZN(n35) );
  AND2_X1 U38 ( .A1(in[12]), .A2(n67), .ZN(n36) );
  AND2_X1 U39 ( .A1(in[13]), .A2(n67), .ZN(n37) );
  AND2_X1 U40 ( .A1(in[14]), .A2(n67), .ZN(n38) );
  AND2_X1 U41 ( .A1(in[15]), .A2(n67), .ZN(n39) );
  AND2_X1 U42 ( .A1(in[16]), .A2(n67), .ZN(n40) );
  AND2_X1 U43 ( .A1(in[17]), .A2(n67), .ZN(n41) );
  AND2_X1 U44 ( .A1(in[18]), .A2(n67), .ZN(n42) );
  AND2_X1 U45 ( .A1(in[19]), .A2(n67), .ZN(n43) );
  AND2_X1 U46 ( .A1(in[20]), .A2(n67), .ZN(n44) );
  AND2_X1 U47 ( .A1(in[21]), .A2(n66), .ZN(n45) );
  AND2_X1 U48 ( .A1(in[22]), .A2(n66), .ZN(n46) );
  AND2_X1 U49 ( .A1(in[23]), .A2(n66), .ZN(n47) );
  AND2_X1 U50 ( .A1(in[24]), .A2(n66), .ZN(n48) );
  AND2_X1 U51 ( .A1(in[25]), .A2(n66), .ZN(n49) );
  AND2_X1 U52 ( .A1(in[26]), .A2(n66), .ZN(n50) );
  AND2_X1 U53 ( .A1(in[27]), .A2(n66), .ZN(n51) );
  AND2_X1 U54 ( .A1(in[28]), .A2(n66), .ZN(n52) );
  AND2_X1 U55 ( .A1(in[29]), .A2(n66), .ZN(n53) );
  AND2_X1 U56 ( .A1(in[30]), .A2(n66), .ZN(n54) );
  AND2_X1 U57 ( .A1(in[31]), .A2(n66), .ZN(n55) );
  AND2_X1 U58 ( .A1(in[0]), .A2(n68), .ZN(n56) );
  AND2_X1 U59 ( .A1(in[1]), .A2(n68), .ZN(n57) );
  AND2_X1 U60 ( .A1(in[2]), .A2(n68), .ZN(n58) );
  AND2_X1 U61 ( .A1(in[3]), .A2(n68), .ZN(n59) );
  AND2_X1 U62 ( .A1(in[4]), .A2(n68), .ZN(n60) );
  AND2_X1 U63 ( .A1(in[5]), .A2(n68), .ZN(n61) );
  AND2_X1 U64 ( .A1(in[6]), .A2(n68), .ZN(n62) );
  AND2_X1 U65 ( .A1(in[7]), .A2(n68), .ZN(n63) );
  AND2_X1 U66 ( .A1(in[8]), .A2(n68), .ZN(n64) );
  AND2_X1 U67 ( .A1(in[9]), .A2(n68), .ZN(n65) );
  BUF_X1 U68 ( .A(n33), .Z(n67) );
  BUF_X1 U69 ( .A(n33), .Z(n66) );
  BUF_X1 U70 ( .A(n33), .Z(n68) );
  INV_X1 U71 ( .A(reset), .ZN(n33) );
endmodule



module BWAdder ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317;
  assign carry[0] = 1'b0;

  XOR2_X1 U256 ( .A(c[9]), .B(n191), .Z(result[9]) );
  XOR2_X1 U257 ( .A(c[8]), .B(n192), .Z(result[8]) );
  XOR2_X1 U258 ( .A(c[7]), .B(n193), .Z(result[7]) );
  XOR2_X1 U259 ( .A(c[6]), .B(n194), .Z(result[6]) );
  XOR2_X1 U260 ( .A(a[63]), .B(n195), .Z(result[63]) );
  XOR2_X1 U261 ( .A(c[63]), .B(b[63]), .Z(n195) );
  XOR2_X1 U262 ( .A(c[62]), .B(n196), .Z(result[62]) );
  XOR2_X1 U263 ( .A(c[61]), .B(n197), .Z(result[61]) );
  XOR2_X1 U264 ( .A(c[60]), .B(n198), .Z(result[60]) );
  XOR2_X1 U265 ( .A(c[5]), .B(n199), .Z(result[5]) );
  XOR2_X1 U266 ( .A(c[59]), .B(n200), .Z(result[59]) );
  XOR2_X1 U267 ( .A(c[58]), .B(n201), .Z(result[58]) );
  XOR2_X1 U268 ( .A(c[57]), .B(n202), .Z(result[57]) );
  XOR2_X1 U269 ( .A(c[56]), .B(n203), .Z(result[56]) );
  XOR2_X1 U270 ( .A(c[55]), .B(n204), .Z(result[55]) );
  XOR2_X1 U271 ( .A(c[54]), .B(n205), .Z(result[54]) );
  XOR2_X1 U272 ( .A(c[53]), .B(n206), .Z(result[53]) );
  XOR2_X1 U273 ( .A(c[52]), .B(n207), .Z(result[52]) );
  XOR2_X1 U274 ( .A(c[51]), .B(n208), .Z(result[51]) );
  XOR2_X1 U275 ( .A(c[50]), .B(n209), .Z(result[50]) );
  XOR2_X1 U276 ( .A(c[4]), .B(n210), .Z(result[4]) );
  XOR2_X1 U277 ( .A(c[49]), .B(n211), .Z(result[49]) );
  XOR2_X1 U278 ( .A(c[48]), .B(n212), .Z(result[48]) );
  XOR2_X1 U279 ( .A(c[47]), .B(n213), .Z(result[47]) );
  XOR2_X1 U280 ( .A(c[46]), .B(n214), .Z(result[46]) );
  XOR2_X1 U281 ( .A(c[45]), .B(n215), .Z(result[45]) );
  XOR2_X1 U282 ( .A(c[44]), .B(n216), .Z(result[44]) );
  XOR2_X1 U283 ( .A(c[43]), .B(n217), .Z(result[43]) );
  XOR2_X1 U284 ( .A(c[42]), .B(n218), .Z(result[42]) );
  XOR2_X1 U285 ( .A(c[41]), .B(n219), .Z(result[41]) );
  XOR2_X1 U286 ( .A(c[40]), .B(n220), .Z(result[40]) );
  XOR2_X1 U287 ( .A(c[3]), .B(n221), .Z(result[3]) );
  XOR2_X1 U288 ( .A(c[39]), .B(n222), .Z(result[39]) );
  XOR2_X1 U289 ( .A(c[38]), .B(n223), .Z(result[38]) );
  XOR2_X1 U290 ( .A(c[37]), .B(n224), .Z(result[37]) );
  XOR2_X1 U291 ( .A(c[36]), .B(n225), .Z(result[36]) );
  XOR2_X1 U292 ( .A(c[35]), .B(n226), .Z(result[35]) );
  XOR2_X1 U293 ( .A(c[34]), .B(n227), .Z(result[34]) );
  XOR2_X1 U294 ( .A(c[33]), .B(n228), .Z(result[33]) );
  XOR2_X1 U295 ( .A(c[32]), .B(n229), .Z(result[32]) );
  XOR2_X1 U296 ( .A(c[31]), .B(n230), .Z(result[31]) );
  XOR2_X1 U297 ( .A(c[30]), .B(n231), .Z(result[30]) );
  XOR2_X1 U298 ( .A(c[2]), .B(n232), .Z(result[2]) );
  XOR2_X1 U299 ( .A(c[29]), .B(n233), .Z(result[29]) );
  XOR2_X1 U300 ( .A(c[28]), .B(n234), .Z(result[28]) );
  XOR2_X1 U301 ( .A(c[27]), .B(n235), .Z(result[27]) );
  XOR2_X1 U302 ( .A(c[26]), .B(n236), .Z(result[26]) );
  XOR2_X1 U303 ( .A(c[25]), .B(n237), .Z(result[25]) );
  XOR2_X1 U304 ( .A(c[24]), .B(n238), .Z(result[24]) );
  XOR2_X1 U305 ( .A(c[23]), .B(n239), .Z(result[23]) );
  XOR2_X1 U306 ( .A(c[22]), .B(n240), .Z(result[22]) );
  XOR2_X1 U307 ( .A(c[21]), .B(n241), .Z(result[21]) );
  XOR2_X1 U308 ( .A(c[20]), .B(n242), .Z(result[20]) );
  XOR2_X1 U309 ( .A(c[1]), .B(n243), .Z(result[1]) );
  XOR2_X1 U310 ( .A(c[19]), .B(n244), .Z(result[19]) );
  XOR2_X1 U311 ( .A(c[18]), .B(n245), .Z(result[18]) );
  XOR2_X1 U312 ( .A(c[17]), .B(n246), .Z(result[17]) );
  XOR2_X1 U313 ( .A(c[16]), .B(n247), .Z(result[16]) );
  XOR2_X1 U314 ( .A(c[15]), .B(n248), .Z(result[15]) );
  XOR2_X1 U315 ( .A(c[14]), .B(n249), .Z(result[14]) );
  XOR2_X1 U316 ( .A(c[13]), .B(n250), .Z(result[13]) );
  XOR2_X1 U317 ( .A(c[12]), .B(n251), .Z(result[12]) );
  XOR2_X1 U318 ( .A(c[11]), .B(n252), .Z(result[11]) );
  XOR2_X1 U319 ( .A(c[10]), .B(n253), .Z(result[10]) );
  XOR2_X1 U320 ( .A(c[0]), .B(n254), .Z(result[0]) );
  INV_X1 U321 ( .A(n255), .ZN(carry[9]) );
  AOI22_X1 U322 ( .A1(b[8]), .A2(a[8]), .B1(n192), .B2(c[8]), .ZN(n255) );
  XOR2_X1 U323 ( .A(a[8]), .B(b[8]), .Z(n192) );
  INV_X1 U324 ( .A(n256), .ZN(carry[8]) );
  AOI22_X1 U325 ( .A1(b[7]), .A2(a[7]), .B1(n193), .B2(c[7]), .ZN(n256) );
  XOR2_X1 U326 ( .A(a[7]), .B(b[7]), .Z(n193) );
  INV_X1 U327 ( .A(n257), .ZN(carry[7]) );
  AOI22_X1 U328 ( .A1(b[6]), .A2(a[6]), .B1(n194), .B2(c[6]), .ZN(n257) );
  XOR2_X1 U329 ( .A(a[6]), .B(b[6]), .Z(n194) );
  INV_X1 U330 ( .A(n258), .ZN(carry[6]) );
  AOI22_X1 U331 ( .A1(b[5]), .A2(a[5]), .B1(n199), .B2(c[5]), .ZN(n258) );
  XOR2_X1 U332 ( .A(a[5]), .B(b[5]), .Z(n199) );
  INV_X1 U333 ( .A(n259), .ZN(carry[63]) );
  AOI22_X1 U334 ( .A1(b[62]), .A2(a[62]), .B1(n196), .B2(c[62]), .ZN(n259) );
  XOR2_X1 U335 ( .A(a[62]), .B(b[62]), .Z(n196) );
  INV_X1 U336 ( .A(n260), .ZN(carry[62]) );
  AOI22_X1 U337 ( .A1(b[61]), .A2(a[61]), .B1(n197), .B2(c[61]), .ZN(n260) );
  XOR2_X1 U338 ( .A(a[61]), .B(b[61]), .Z(n197) );
  INV_X1 U339 ( .A(n261), .ZN(carry[61]) );
  AOI22_X1 U340 ( .A1(b[60]), .A2(a[60]), .B1(n198), .B2(c[60]), .ZN(n261) );
  XOR2_X1 U341 ( .A(a[60]), .B(b[60]), .Z(n198) );
  INV_X1 U342 ( .A(n262), .ZN(carry[60]) );
  AOI22_X1 U343 ( .A1(b[59]), .A2(a[59]), .B1(n200), .B2(c[59]), .ZN(n262) );
  XOR2_X1 U344 ( .A(a[59]), .B(b[59]), .Z(n200) );
  INV_X1 U345 ( .A(n263), .ZN(carry[5]) );
  AOI22_X1 U346 ( .A1(b[4]), .A2(a[4]), .B1(n210), .B2(c[4]), .ZN(n263) );
  XOR2_X1 U347 ( .A(a[4]), .B(b[4]), .Z(n210) );
  INV_X1 U348 ( .A(n264), .ZN(carry[59]) );
  AOI22_X1 U349 ( .A1(b[58]), .A2(a[58]), .B1(n201), .B2(c[58]), .ZN(n264) );
  XOR2_X1 U350 ( .A(a[58]), .B(b[58]), .Z(n201) );
  INV_X1 U351 ( .A(n265), .ZN(carry[58]) );
  AOI22_X1 U352 ( .A1(b[57]), .A2(a[57]), .B1(n202), .B2(c[57]), .ZN(n265) );
  XOR2_X1 U353 ( .A(a[57]), .B(b[57]), .Z(n202) );
  INV_X1 U354 ( .A(n266), .ZN(carry[57]) );
  AOI22_X1 U355 ( .A1(b[56]), .A2(a[56]), .B1(n203), .B2(c[56]), .ZN(n266) );
  XOR2_X1 U356 ( .A(a[56]), .B(b[56]), .Z(n203) );
  INV_X1 U357 ( .A(n267), .ZN(carry[56]) );
  AOI22_X1 U358 ( .A1(b[55]), .A2(a[55]), .B1(n204), .B2(c[55]), .ZN(n267) );
  XOR2_X1 U359 ( .A(a[55]), .B(b[55]), .Z(n204) );
  INV_X1 U360 ( .A(n268), .ZN(carry[55]) );
  AOI22_X1 U361 ( .A1(b[54]), .A2(a[54]), .B1(n205), .B2(c[54]), .ZN(n268) );
  XOR2_X1 U362 ( .A(a[54]), .B(b[54]), .Z(n205) );
  INV_X1 U363 ( .A(n269), .ZN(carry[54]) );
  AOI22_X1 U364 ( .A1(b[53]), .A2(a[53]), .B1(n206), .B2(c[53]), .ZN(n269) );
  XOR2_X1 U365 ( .A(a[53]), .B(b[53]), .Z(n206) );
  INV_X1 U366 ( .A(n270), .ZN(carry[53]) );
  AOI22_X1 U367 ( .A1(b[52]), .A2(a[52]), .B1(n207), .B2(c[52]), .ZN(n270) );
  XOR2_X1 U368 ( .A(a[52]), .B(b[52]), .Z(n207) );
  INV_X1 U369 ( .A(n271), .ZN(carry[52]) );
  AOI22_X1 U370 ( .A1(b[51]), .A2(a[51]), .B1(n208), .B2(c[51]), .ZN(n271) );
  XOR2_X1 U371 ( .A(a[51]), .B(b[51]), .Z(n208) );
  INV_X1 U372 ( .A(n272), .ZN(carry[51]) );
  AOI22_X1 U373 ( .A1(b[50]), .A2(a[50]), .B1(n209), .B2(c[50]), .ZN(n272) );
  XOR2_X1 U374 ( .A(a[50]), .B(b[50]), .Z(n209) );
  INV_X1 U375 ( .A(n273), .ZN(carry[50]) );
  AOI22_X1 U376 ( .A1(b[49]), .A2(a[49]), .B1(n211), .B2(c[49]), .ZN(n273) );
  XOR2_X1 U377 ( .A(a[49]), .B(b[49]), .Z(n211) );
  INV_X1 U378 ( .A(n274), .ZN(carry[4]) );
  AOI22_X1 U379 ( .A1(b[3]), .A2(a[3]), .B1(n221), .B2(c[3]), .ZN(n274) );
  XOR2_X1 U380 ( .A(a[3]), .B(b[3]), .Z(n221) );
  INV_X1 U381 ( .A(n275), .ZN(carry[49]) );
  AOI22_X1 U382 ( .A1(b[48]), .A2(a[48]), .B1(n212), .B2(c[48]), .ZN(n275) );
  XOR2_X1 U383 ( .A(a[48]), .B(b[48]), .Z(n212) );
  INV_X1 U384 ( .A(n276), .ZN(carry[48]) );
  AOI22_X1 U385 ( .A1(b[47]), .A2(a[47]), .B1(n213), .B2(c[47]), .ZN(n276) );
  XOR2_X1 U386 ( .A(a[47]), .B(b[47]), .Z(n213) );
  INV_X1 U387 ( .A(n277), .ZN(carry[47]) );
  AOI22_X1 U388 ( .A1(b[46]), .A2(a[46]), .B1(n214), .B2(c[46]), .ZN(n277) );
  XOR2_X1 U389 ( .A(a[46]), .B(b[46]), .Z(n214) );
  INV_X1 U390 ( .A(n278), .ZN(carry[46]) );
  AOI22_X1 U391 ( .A1(b[45]), .A2(a[45]), .B1(n215), .B2(c[45]), .ZN(n278) );
  XOR2_X1 U392 ( .A(a[45]), .B(b[45]), .Z(n215) );
  INV_X1 U393 ( .A(n279), .ZN(carry[45]) );
  AOI22_X1 U394 ( .A1(b[44]), .A2(a[44]), .B1(n216), .B2(c[44]), .ZN(n279) );
  XOR2_X1 U395 ( .A(a[44]), .B(b[44]), .Z(n216) );
  INV_X1 U396 ( .A(n280), .ZN(carry[44]) );
  AOI22_X1 U397 ( .A1(b[43]), .A2(a[43]), .B1(n217), .B2(c[43]), .ZN(n280) );
  XOR2_X1 U398 ( .A(a[43]), .B(b[43]), .Z(n217) );
  INV_X1 U399 ( .A(n281), .ZN(carry[43]) );
  AOI22_X1 U400 ( .A1(b[42]), .A2(a[42]), .B1(n218), .B2(c[42]), .ZN(n281) );
  XOR2_X1 U401 ( .A(a[42]), .B(b[42]), .Z(n218) );
  INV_X1 U402 ( .A(n282), .ZN(carry[42]) );
  AOI22_X1 U403 ( .A1(b[41]), .A2(a[41]), .B1(n219), .B2(c[41]), .ZN(n282) );
  XOR2_X1 U404 ( .A(a[41]), .B(b[41]), .Z(n219) );
  INV_X1 U405 ( .A(n283), .ZN(carry[41]) );
  AOI22_X1 U406 ( .A1(b[40]), .A2(a[40]), .B1(n220), .B2(c[40]), .ZN(n283) );
  XOR2_X1 U407 ( .A(a[40]), .B(b[40]), .Z(n220) );
  INV_X1 U408 ( .A(n284), .ZN(carry[40]) );
  AOI22_X1 U409 ( .A1(b[39]), .A2(a[39]), .B1(n222), .B2(c[39]), .ZN(n284) );
  XOR2_X1 U410 ( .A(a[39]), .B(b[39]), .Z(n222) );
  INV_X1 U411 ( .A(n285), .ZN(carry[3]) );
  AOI22_X1 U412 ( .A1(b[2]), .A2(a[2]), .B1(n232), .B2(c[2]), .ZN(n285) );
  XOR2_X1 U413 ( .A(a[2]), .B(b[2]), .Z(n232) );
  INV_X1 U414 ( .A(n286), .ZN(carry[39]) );
  AOI22_X1 U415 ( .A1(b[38]), .A2(a[38]), .B1(n223), .B2(c[38]), .ZN(n286) );
  XOR2_X1 U416 ( .A(a[38]), .B(b[38]), .Z(n223) );
  INV_X1 U417 ( .A(n287), .ZN(carry[38]) );
  AOI22_X1 U418 ( .A1(b[37]), .A2(a[37]), .B1(n224), .B2(c[37]), .ZN(n287) );
  XOR2_X1 U419 ( .A(a[37]), .B(b[37]), .Z(n224) );
  INV_X1 U420 ( .A(n288), .ZN(carry[37]) );
  AOI22_X1 U421 ( .A1(b[36]), .A2(a[36]), .B1(n225), .B2(c[36]), .ZN(n288) );
  XOR2_X1 U422 ( .A(a[36]), .B(b[36]), .Z(n225) );
  INV_X1 U423 ( .A(n289), .ZN(carry[36]) );
  AOI22_X1 U424 ( .A1(b[35]), .A2(a[35]), .B1(n226), .B2(c[35]), .ZN(n289) );
  XOR2_X1 U425 ( .A(a[35]), .B(b[35]), .Z(n226) );
  INV_X1 U426 ( .A(n290), .ZN(carry[35]) );
  AOI22_X1 U427 ( .A1(b[34]), .A2(a[34]), .B1(n227), .B2(c[34]), .ZN(n290) );
  XOR2_X1 U428 ( .A(a[34]), .B(b[34]), .Z(n227) );
  INV_X1 U429 ( .A(n291), .ZN(carry[34]) );
  AOI22_X1 U430 ( .A1(b[33]), .A2(a[33]), .B1(n228), .B2(c[33]), .ZN(n291) );
  XOR2_X1 U431 ( .A(a[33]), .B(b[33]), .Z(n228) );
  INV_X1 U432 ( .A(n292), .ZN(carry[33]) );
  AOI22_X1 U433 ( .A1(b[32]), .A2(a[32]), .B1(n229), .B2(c[32]), .ZN(n292) );
  XOR2_X1 U434 ( .A(a[32]), .B(b[32]), .Z(n229) );
  INV_X1 U435 ( .A(n293), .ZN(carry[32]) );
  AOI22_X1 U436 ( .A1(b[31]), .A2(a[31]), .B1(n230), .B2(c[31]), .ZN(n293) );
  XOR2_X1 U437 ( .A(a[31]), .B(b[31]), .Z(n230) );
  INV_X1 U438 ( .A(n294), .ZN(carry[31]) );
  AOI22_X1 U439 ( .A1(b[30]), .A2(a[30]), .B1(n231), .B2(c[30]), .ZN(n294) );
  XOR2_X1 U440 ( .A(a[30]), .B(b[30]), .Z(n231) );
  INV_X1 U441 ( .A(n295), .ZN(carry[30]) );
  AOI22_X1 U442 ( .A1(b[29]), .A2(a[29]), .B1(n233), .B2(c[29]), .ZN(n295) );
  XOR2_X1 U443 ( .A(a[29]), .B(b[29]), .Z(n233) );
  INV_X1 U444 ( .A(n296), .ZN(carry[2]) );
  AOI22_X1 U445 ( .A1(b[1]), .A2(a[1]), .B1(n243), .B2(c[1]), .ZN(n296) );
  XOR2_X1 U446 ( .A(a[1]), .B(b[1]), .Z(n243) );
  INV_X1 U447 ( .A(n297), .ZN(carry[29]) );
  AOI22_X1 U448 ( .A1(b[28]), .A2(a[28]), .B1(n234), .B2(c[28]), .ZN(n297) );
  XOR2_X1 U449 ( .A(a[28]), .B(b[28]), .Z(n234) );
  INV_X1 U450 ( .A(n298), .ZN(carry[28]) );
  AOI22_X1 U451 ( .A1(b[27]), .A2(a[27]), .B1(n235), .B2(c[27]), .ZN(n298) );
  XOR2_X1 U452 ( .A(a[27]), .B(b[27]), .Z(n235) );
  INV_X1 U453 ( .A(n299), .ZN(carry[27]) );
  AOI22_X1 U454 ( .A1(b[26]), .A2(a[26]), .B1(n236), .B2(c[26]), .ZN(n299) );
  XOR2_X1 U455 ( .A(a[26]), .B(b[26]), .Z(n236) );
  INV_X1 U456 ( .A(n300), .ZN(carry[26]) );
  AOI22_X1 U457 ( .A1(b[25]), .A2(a[25]), .B1(n237), .B2(c[25]), .ZN(n300) );
  XOR2_X1 U458 ( .A(a[25]), .B(b[25]), .Z(n237) );
  INV_X1 U459 ( .A(n301), .ZN(carry[25]) );
  AOI22_X1 U460 ( .A1(b[24]), .A2(a[24]), .B1(n238), .B2(c[24]), .ZN(n301) );
  XOR2_X1 U461 ( .A(a[24]), .B(b[24]), .Z(n238) );
  INV_X1 U462 ( .A(n302), .ZN(carry[24]) );
  AOI22_X1 U463 ( .A1(b[23]), .A2(a[23]), .B1(n239), .B2(c[23]), .ZN(n302) );
  XOR2_X1 U464 ( .A(a[23]), .B(b[23]), .Z(n239) );
  INV_X1 U465 ( .A(n303), .ZN(carry[23]) );
  AOI22_X1 U466 ( .A1(b[22]), .A2(a[22]), .B1(n240), .B2(c[22]), .ZN(n303) );
  XOR2_X1 U467 ( .A(a[22]), .B(b[22]), .Z(n240) );
  INV_X1 U468 ( .A(n304), .ZN(carry[22]) );
  AOI22_X1 U469 ( .A1(b[21]), .A2(a[21]), .B1(n241), .B2(c[21]), .ZN(n304) );
  XOR2_X1 U470 ( .A(a[21]), .B(b[21]), .Z(n241) );
  INV_X1 U471 ( .A(n305), .ZN(carry[21]) );
  AOI22_X1 U472 ( .A1(b[20]), .A2(a[20]), .B1(n242), .B2(c[20]), .ZN(n305) );
  XOR2_X1 U473 ( .A(a[20]), .B(b[20]), .Z(n242) );
  INV_X1 U474 ( .A(n306), .ZN(carry[20]) );
  AOI22_X1 U475 ( .A1(b[19]), .A2(a[19]), .B1(n244), .B2(c[19]), .ZN(n306) );
  XOR2_X1 U476 ( .A(a[19]), .B(b[19]), .Z(n244) );
  INV_X1 U477 ( .A(n307), .ZN(carry[1]) );
  AOI22_X1 U478 ( .A1(b[0]), .A2(a[0]), .B1(n254), .B2(c[0]), .ZN(n307) );
  XOR2_X1 U479 ( .A(a[0]), .B(b[0]), .Z(n254) );
  INV_X1 U480 ( .A(n308), .ZN(carry[19]) );
  AOI22_X1 U481 ( .A1(b[18]), .A2(a[18]), .B1(n245), .B2(c[18]), .ZN(n308) );
  XOR2_X1 U482 ( .A(a[18]), .B(b[18]), .Z(n245) );
  INV_X1 U483 ( .A(n309), .ZN(carry[18]) );
  AOI22_X1 U484 ( .A1(b[17]), .A2(a[17]), .B1(n246), .B2(c[17]), .ZN(n309) );
  XOR2_X1 U485 ( .A(a[17]), .B(b[17]), .Z(n246) );
  INV_X1 U486 ( .A(n310), .ZN(carry[17]) );
  AOI22_X1 U487 ( .A1(b[16]), .A2(a[16]), .B1(n247), .B2(c[16]), .ZN(n310) );
  XOR2_X1 U488 ( .A(a[16]), .B(b[16]), .Z(n247) );
  INV_X1 U489 ( .A(n311), .ZN(carry[16]) );
  AOI22_X1 U490 ( .A1(b[15]), .A2(a[15]), .B1(n248), .B2(c[15]), .ZN(n311) );
  XOR2_X1 U491 ( .A(a[15]), .B(b[15]), .Z(n248) );
  INV_X1 U492 ( .A(n312), .ZN(carry[15]) );
  AOI22_X1 U493 ( .A1(b[14]), .A2(a[14]), .B1(n249), .B2(c[14]), .ZN(n312) );
  XOR2_X1 U494 ( .A(a[14]), .B(b[14]), .Z(n249) );
  INV_X1 U495 ( .A(n313), .ZN(carry[14]) );
  AOI22_X1 U496 ( .A1(b[13]), .A2(a[13]), .B1(n250), .B2(c[13]), .ZN(n313) );
  XOR2_X1 U497 ( .A(a[13]), .B(b[13]), .Z(n250) );
  INV_X1 U498 ( .A(n314), .ZN(carry[13]) );
  AOI22_X1 U499 ( .A1(b[12]), .A2(a[12]), .B1(n251), .B2(c[12]), .ZN(n314) );
  XOR2_X1 U500 ( .A(a[12]), .B(b[12]), .Z(n251) );
  INV_X1 U501 ( .A(n315), .ZN(carry[12]) );
  AOI22_X1 U502 ( .A1(b[11]), .A2(a[11]), .B1(n252), .B2(c[11]), .ZN(n315) );
  XOR2_X1 U503 ( .A(a[11]), .B(b[11]), .Z(n252) );
  INV_X1 U504 ( .A(n316), .ZN(carry[11]) );
  AOI22_X1 U505 ( .A1(b[10]), .A2(a[10]), .B1(n253), .B2(c[10]), .ZN(n316) );
  XOR2_X1 U506 ( .A(a[10]), .B(b[10]), .Z(n253) );
  INV_X1 U507 ( .A(n317), .ZN(carry[10]) );
  AOI22_X1 U508 ( .A1(b[9]), .A2(a[9]), .B1(n191), .B2(c[9]), .ZN(n317) );
  XOR2_X1 U509 ( .A(a[9]), .B(b[9]), .Z(n191) );
endmodule


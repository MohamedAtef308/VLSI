
module BWAdder_0 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module FullAdder_0 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_3 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_4 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_5 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_6 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_7 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_8 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_9 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_10 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_11 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_12 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_13 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_14 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_15 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_16 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_17 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_18 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_19 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_20 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_21 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_22 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_23 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_24 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_25 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_26 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_27 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_28 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_29 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_30 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_31 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_32 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_33 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_34 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_35 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_36 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_37 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_38 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_39 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_40 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_41 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_42 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_43 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_44 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_45 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_46 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_47 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_48 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_49 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_50 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_51 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_52 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_53 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_54 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_55 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_56 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_57 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_58 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_59 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_60 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_61 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_62 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_63 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_64 ( a, b, cin, sum, cout, overflow );
  input [63:0] a;
  input [63:0] b;
  output [63:0] sum;
  input cin;
  output cout, overflow;
  wire   n1, n2;
  wire   [62:0] passCout;

  FullAdder_0 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_63 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_62 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_61 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_60 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_59 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_58 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_57 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_56 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_55 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_54 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_53 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_52 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_51 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_50 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_49 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_48 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_47 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_46 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_45 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_44 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_43 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_42 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_41 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_40 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_39 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_38 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_37 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_36 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_35 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_34 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_33 bit_gen_31__bit ( .a(a[31]), .b(b[31]), .cin(passCout[30]), 
        .sum(sum[31]), .cout(passCout[31]) );
  FullAdder_32 bit_gen_32__bit ( .a(a[32]), .b(b[32]), .cin(passCout[31]), 
        .sum(sum[32]), .cout(passCout[32]) );
  FullAdder_31 bit_gen_33__bit ( .a(a[33]), .b(b[33]), .cin(passCout[32]), 
        .sum(sum[33]), .cout(passCout[33]) );
  FullAdder_30 bit_gen_34__bit ( .a(a[34]), .b(b[34]), .cin(passCout[33]), 
        .sum(sum[34]), .cout(passCout[34]) );
  FullAdder_29 bit_gen_35__bit ( .a(a[35]), .b(b[35]), .cin(passCout[34]), 
        .sum(sum[35]), .cout(passCout[35]) );
  FullAdder_28 bit_gen_36__bit ( .a(a[36]), .b(b[36]), .cin(passCout[35]), 
        .sum(sum[36]), .cout(passCout[36]) );
  FullAdder_27 bit_gen_37__bit ( .a(a[37]), .b(b[37]), .cin(passCout[36]), 
        .sum(sum[37]), .cout(passCout[37]) );
  FullAdder_26 bit_gen_38__bit ( .a(a[38]), .b(b[38]), .cin(passCout[37]), 
        .sum(sum[38]), .cout(passCout[38]) );
  FullAdder_25 bit_gen_39__bit ( .a(a[39]), .b(b[39]), .cin(passCout[38]), 
        .sum(sum[39]), .cout(passCout[39]) );
  FullAdder_24 bit_gen_40__bit ( .a(a[40]), .b(b[40]), .cin(passCout[39]), 
        .sum(sum[40]), .cout(passCout[40]) );
  FullAdder_23 bit_gen_41__bit ( .a(a[41]), .b(b[41]), .cin(passCout[40]), 
        .sum(sum[41]), .cout(passCout[41]) );
  FullAdder_22 bit_gen_42__bit ( .a(a[42]), .b(b[42]), .cin(passCout[41]), 
        .sum(sum[42]), .cout(passCout[42]) );
  FullAdder_21 bit_gen_43__bit ( .a(a[43]), .b(b[43]), .cin(passCout[42]), 
        .sum(sum[43]), .cout(passCout[43]) );
  FullAdder_20 bit_gen_44__bit ( .a(a[44]), .b(b[44]), .cin(passCout[43]), 
        .sum(sum[44]), .cout(passCout[44]) );
  FullAdder_19 bit_gen_45__bit ( .a(a[45]), .b(b[45]), .cin(passCout[44]), 
        .sum(sum[45]), .cout(passCout[45]) );
  FullAdder_18 bit_gen_46__bit ( .a(a[46]), .b(b[46]), .cin(passCout[45]), 
        .sum(sum[46]), .cout(passCout[46]) );
  FullAdder_17 bit_gen_47__bit ( .a(a[47]), .b(b[47]), .cin(passCout[46]), 
        .sum(sum[47]), .cout(passCout[47]) );
  FullAdder_16 bit_gen_48__bit ( .a(a[48]), .b(b[48]), .cin(passCout[47]), 
        .sum(sum[48]), .cout(passCout[48]) );
  FullAdder_15 bit_gen_49__bit ( .a(a[49]), .b(b[49]), .cin(passCout[48]), 
        .sum(sum[49]), .cout(passCout[49]) );
  FullAdder_14 bit_gen_50__bit ( .a(a[50]), .b(b[50]), .cin(passCout[49]), 
        .sum(sum[50]), .cout(passCout[50]) );
  FullAdder_13 bit_gen_51__bit ( .a(a[51]), .b(b[51]), .cin(passCout[50]), 
        .sum(sum[51]), .cout(passCout[51]) );
  FullAdder_12 bit_gen_52__bit ( .a(a[52]), .b(b[52]), .cin(passCout[51]), 
        .sum(sum[52]), .cout(passCout[52]) );
  FullAdder_11 bit_gen_53__bit ( .a(a[53]), .b(b[53]), .cin(passCout[52]), 
        .sum(sum[53]), .cout(passCout[53]) );
  FullAdder_10 bit_gen_54__bit ( .a(a[54]), .b(b[54]), .cin(passCout[53]), 
        .sum(sum[54]), .cout(passCout[54]) );
  FullAdder_9 bit_gen_55__bit ( .a(a[55]), .b(b[55]), .cin(passCout[54]), 
        .sum(sum[55]), .cout(passCout[55]) );
  FullAdder_8 bit_gen_56__bit ( .a(a[56]), .b(b[56]), .cin(passCout[55]), 
        .sum(sum[56]), .cout(passCout[56]) );
  FullAdder_7 bit_gen_57__bit ( .a(a[57]), .b(b[57]), .cin(passCout[56]), 
        .sum(sum[57]), .cout(passCout[57]) );
  FullAdder_6 bit_gen_58__bit ( .a(a[58]), .b(b[58]), .cin(passCout[57]), 
        .sum(sum[58]), .cout(passCout[58]) );
  FullAdder_5 bit_gen_59__bit ( .a(a[59]), .b(b[59]), .cin(passCout[58]), 
        .sum(sum[59]), .cout(passCout[59]) );
  FullAdder_4 bit_gen_60__bit ( .a(a[60]), .b(b[60]), .cin(passCout[59]), 
        .sum(sum[60]), .cout(passCout[60]) );
  FullAdder_3 bit_gen_61__bit ( .a(a[61]), .b(b[61]), .cin(passCout[60]), 
        .sum(sum[61]), .cout(passCout[61]) );
  FullAdder_2 bit_gen_62__bit ( .a(a[62]), .b(b[62]), .cin(passCout[61]), 
        .sum(sum[62]), .cout(passCout[62]) );
  FullAdder_1 bit63 ( .a(a[63]), .b(b[63]), .cin(passCout[62]), .sum(sum[63]), 
        .cout(cout) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(overflow) );
  XOR2_X1 U2 ( .A(b[63]), .B(a[63]), .Z(n2) );
  XNOR2_X1 U3 ( .A(a[63]), .B(sum[63]), .ZN(n1) );
endmodule


module BWAdder_1 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_2 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_3 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_4 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_5 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_6 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_7 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_8 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_9 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_10 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_11 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_12 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_13 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_14 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_15 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_16 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_17 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_18 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_19 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_20 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_21 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_22 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_23 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_24 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_25 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_26 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_27 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_28 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_29 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_30 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_31 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_32 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_33 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_34 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_35 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_36 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_37 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_38 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_39 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_40 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_41 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_42 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_43 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_44 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_45 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_46 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_47 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_48 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_49 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_50 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_51 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_52 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_53 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_54 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_55 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_56 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_57 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_58 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_59 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_60 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module BWAdder_61 ( a, b, c, result, carry );
  input [63:0] a;
  input [63:0] b;
  input [63:0] c;
  output [63:0] result;
  output [63:0] carry;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127;
  assign carry[0] = 1'b0;

  XOR2_X1 U2 ( .A(c[9]), .B(n1), .Z(result[9]) );
  XOR2_X1 U3 ( .A(c[8]), .B(n2), .Z(result[8]) );
  XOR2_X1 U4 ( .A(c[7]), .B(n3), .Z(result[7]) );
  XOR2_X1 U5 ( .A(c[6]), .B(n4), .Z(result[6]) );
  XOR2_X1 U6 ( .A(a[63]), .B(n5), .Z(result[63]) );
  XOR2_X1 U7 ( .A(c[63]), .B(b[63]), .Z(n5) );
  XOR2_X1 U8 ( .A(c[62]), .B(n6), .Z(result[62]) );
  XOR2_X1 U9 ( .A(c[61]), .B(n7), .Z(result[61]) );
  XOR2_X1 U10 ( .A(c[60]), .B(n8), .Z(result[60]) );
  XOR2_X1 U11 ( .A(c[5]), .B(n9), .Z(result[5]) );
  XOR2_X1 U12 ( .A(c[59]), .B(n10), .Z(result[59]) );
  XOR2_X1 U13 ( .A(c[58]), .B(n11), .Z(result[58]) );
  XOR2_X1 U14 ( .A(c[57]), .B(n12), .Z(result[57]) );
  XOR2_X1 U15 ( .A(c[56]), .B(n13), .Z(result[56]) );
  XOR2_X1 U16 ( .A(c[55]), .B(n14), .Z(result[55]) );
  XOR2_X1 U17 ( .A(c[54]), .B(n15), .Z(result[54]) );
  XOR2_X1 U18 ( .A(c[53]), .B(n16), .Z(result[53]) );
  XOR2_X1 U19 ( .A(c[52]), .B(n17), .Z(result[52]) );
  XOR2_X1 U20 ( .A(c[51]), .B(n18), .Z(result[51]) );
  XOR2_X1 U21 ( .A(c[50]), .B(n19), .Z(result[50]) );
  XOR2_X1 U22 ( .A(c[4]), .B(n20), .Z(result[4]) );
  XOR2_X1 U23 ( .A(c[49]), .B(n21), .Z(result[49]) );
  XOR2_X1 U24 ( .A(c[48]), .B(n22), .Z(result[48]) );
  XOR2_X1 U25 ( .A(c[47]), .B(n23), .Z(result[47]) );
  XOR2_X1 U26 ( .A(c[46]), .B(n24), .Z(result[46]) );
  XOR2_X1 U27 ( .A(c[45]), .B(n25), .Z(result[45]) );
  XOR2_X1 U28 ( .A(c[44]), .B(n26), .Z(result[44]) );
  XOR2_X1 U29 ( .A(c[43]), .B(n27), .Z(result[43]) );
  XOR2_X1 U30 ( .A(c[42]), .B(n28), .Z(result[42]) );
  XOR2_X1 U31 ( .A(c[41]), .B(n29), .Z(result[41]) );
  XOR2_X1 U32 ( .A(c[40]), .B(n30), .Z(result[40]) );
  XOR2_X1 U33 ( .A(c[3]), .B(n31), .Z(result[3]) );
  XOR2_X1 U34 ( .A(c[39]), .B(n32), .Z(result[39]) );
  XOR2_X1 U35 ( .A(c[38]), .B(n33), .Z(result[38]) );
  XOR2_X1 U36 ( .A(c[37]), .B(n34), .Z(result[37]) );
  XOR2_X1 U37 ( .A(c[36]), .B(n35), .Z(result[36]) );
  XOR2_X1 U38 ( .A(c[35]), .B(n36), .Z(result[35]) );
  XOR2_X1 U39 ( .A(c[34]), .B(n37), .Z(result[34]) );
  XOR2_X1 U40 ( .A(c[33]), .B(n38), .Z(result[33]) );
  XOR2_X1 U41 ( .A(c[32]), .B(n39), .Z(result[32]) );
  XOR2_X1 U42 ( .A(c[31]), .B(n40), .Z(result[31]) );
  XOR2_X1 U43 ( .A(c[30]), .B(n41), .Z(result[30]) );
  XOR2_X1 U44 ( .A(c[2]), .B(n42), .Z(result[2]) );
  XOR2_X1 U45 ( .A(c[29]), .B(n43), .Z(result[29]) );
  XOR2_X1 U46 ( .A(c[28]), .B(n44), .Z(result[28]) );
  XOR2_X1 U47 ( .A(c[27]), .B(n45), .Z(result[27]) );
  XOR2_X1 U48 ( .A(c[26]), .B(n46), .Z(result[26]) );
  XOR2_X1 U49 ( .A(c[25]), .B(n47), .Z(result[25]) );
  XOR2_X1 U50 ( .A(c[24]), .B(n48), .Z(result[24]) );
  XOR2_X1 U51 ( .A(c[23]), .B(n49), .Z(result[23]) );
  XOR2_X1 U52 ( .A(c[22]), .B(n50), .Z(result[22]) );
  XOR2_X1 U53 ( .A(c[21]), .B(n51), .Z(result[21]) );
  XOR2_X1 U54 ( .A(c[20]), .B(n52), .Z(result[20]) );
  XOR2_X1 U55 ( .A(c[1]), .B(n53), .Z(result[1]) );
  XOR2_X1 U56 ( .A(c[19]), .B(n54), .Z(result[19]) );
  XOR2_X1 U57 ( .A(c[18]), .B(n55), .Z(result[18]) );
  XOR2_X1 U58 ( .A(c[17]), .B(n56), .Z(result[17]) );
  XOR2_X1 U59 ( .A(c[16]), .B(n57), .Z(result[16]) );
  XOR2_X1 U60 ( .A(c[15]), .B(n58), .Z(result[15]) );
  XOR2_X1 U61 ( .A(c[14]), .B(n59), .Z(result[14]) );
  XOR2_X1 U62 ( .A(c[13]), .B(n60), .Z(result[13]) );
  XOR2_X1 U63 ( .A(c[12]), .B(n61), .Z(result[12]) );
  XOR2_X1 U64 ( .A(c[11]), .B(n62), .Z(result[11]) );
  XOR2_X1 U65 ( .A(c[10]), .B(n63), .Z(result[10]) );
  XOR2_X1 U66 ( .A(c[0]), .B(n64), .Z(result[0]) );
  INV_X1 U67 ( .A(n65), .ZN(carry[9]) );
  AOI22_X1 U68 ( .A1(b[8]), .A2(a[8]), .B1(n2), .B2(c[8]), .ZN(n65) );
  XOR2_X1 U69 ( .A(a[8]), .B(b[8]), .Z(n2) );
  INV_X1 U70 ( .A(n66), .ZN(carry[8]) );
  AOI22_X1 U71 ( .A1(b[7]), .A2(a[7]), .B1(n3), .B2(c[7]), .ZN(n66) );
  XOR2_X1 U72 ( .A(a[7]), .B(b[7]), .Z(n3) );
  INV_X1 U73 ( .A(n67), .ZN(carry[7]) );
  AOI22_X1 U74 ( .A1(b[6]), .A2(a[6]), .B1(n4), .B2(c[6]), .ZN(n67) );
  XOR2_X1 U75 ( .A(a[6]), .B(b[6]), .Z(n4) );
  INV_X1 U76 ( .A(n68), .ZN(carry[6]) );
  AOI22_X1 U77 ( .A1(b[5]), .A2(a[5]), .B1(n9), .B2(c[5]), .ZN(n68) );
  XOR2_X1 U78 ( .A(a[5]), .B(b[5]), .Z(n9) );
  INV_X1 U79 ( .A(n69), .ZN(carry[63]) );
  AOI22_X1 U80 ( .A1(b[62]), .A2(a[62]), .B1(n6), .B2(c[62]), .ZN(n69) );
  XOR2_X1 U81 ( .A(a[62]), .B(b[62]), .Z(n6) );
  INV_X1 U82 ( .A(n70), .ZN(carry[62]) );
  AOI22_X1 U83 ( .A1(b[61]), .A2(a[61]), .B1(n7), .B2(c[61]), .ZN(n70) );
  XOR2_X1 U84 ( .A(a[61]), .B(b[61]), .Z(n7) );
  INV_X1 U85 ( .A(n71), .ZN(carry[61]) );
  AOI22_X1 U86 ( .A1(b[60]), .A2(a[60]), .B1(n8), .B2(c[60]), .ZN(n71) );
  XOR2_X1 U87 ( .A(a[60]), .B(b[60]), .Z(n8) );
  INV_X1 U88 ( .A(n72), .ZN(carry[60]) );
  AOI22_X1 U89 ( .A1(b[59]), .A2(a[59]), .B1(n10), .B2(c[59]), .ZN(n72) );
  XOR2_X1 U90 ( .A(a[59]), .B(b[59]), .Z(n10) );
  INV_X1 U91 ( .A(n73), .ZN(carry[5]) );
  AOI22_X1 U92 ( .A1(b[4]), .A2(a[4]), .B1(n20), .B2(c[4]), .ZN(n73) );
  XOR2_X1 U93 ( .A(a[4]), .B(b[4]), .Z(n20) );
  INV_X1 U94 ( .A(n74), .ZN(carry[59]) );
  AOI22_X1 U95 ( .A1(b[58]), .A2(a[58]), .B1(n11), .B2(c[58]), .ZN(n74) );
  XOR2_X1 U96 ( .A(a[58]), .B(b[58]), .Z(n11) );
  INV_X1 U97 ( .A(n75), .ZN(carry[58]) );
  AOI22_X1 U98 ( .A1(b[57]), .A2(a[57]), .B1(n12), .B2(c[57]), .ZN(n75) );
  XOR2_X1 U99 ( .A(a[57]), .B(b[57]), .Z(n12) );
  INV_X1 U100 ( .A(n76), .ZN(carry[57]) );
  AOI22_X1 U101 ( .A1(b[56]), .A2(a[56]), .B1(n13), .B2(c[56]), .ZN(n76) );
  XOR2_X1 U102 ( .A(a[56]), .B(b[56]), .Z(n13) );
  INV_X1 U103 ( .A(n77), .ZN(carry[56]) );
  AOI22_X1 U104 ( .A1(b[55]), .A2(a[55]), .B1(n14), .B2(c[55]), .ZN(n77) );
  XOR2_X1 U105 ( .A(a[55]), .B(b[55]), .Z(n14) );
  INV_X1 U106 ( .A(n78), .ZN(carry[55]) );
  AOI22_X1 U107 ( .A1(b[54]), .A2(a[54]), .B1(n15), .B2(c[54]), .ZN(n78) );
  XOR2_X1 U108 ( .A(a[54]), .B(b[54]), .Z(n15) );
  INV_X1 U109 ( .A(n79), .ZN(carry[54]) );
  AOI22_X1 U110 ( .A1(b[53]), .A2(a[53]), .B1(n16), .B2(c[53]), .ZN(n79) );
  XOR2_X1 U111 ( .A(a[53]), .B(b[53]), .Z(n16) );
  INV_X1 U112 ( .A(n80), .ZN(carry[53]) );
  AOI22_X1 U113 ( .A1(b[52]), .A2(a[52]), .B1(n17), .B2(c[52]), .ZN(n80) );
  XOR2_X1 U114 ( .A(a[52]), .B(b[52]), .Z(n17) );
  INV_X1 U115 ( .A(n81), .ZN(carry[52]) );
  AOI22_X1 U116 ( .A1(b[51]), .A2(a[51]), .B1(n18), .B2(c[51]), .ZN(n81) );
  XOR2_X1 U117 ( .A(a[51]), .B(b[51]), .Z(n18) );
  INV_X1 U118 ( .A(n82), .ZN(carry[51]) );
  AOI22_X1 U119 ( .A1(b[50]), .A2(a[50]), .B1(n19), .B2(c[50]), .ZN(n82) );
  XOR2_X1 U120 ( .A(a[50]), .B(b[50]), .Z(n19) );
  INV_X1 U121 ( .A(n83), .ZN(carry[50]) );
  AOI22_X1 U122 ( .A1(b[49]), .A2(a[49]), .B1(n21), .B2(c[49]), .ZN(n83) );
  XOR2_X1 U123 ( .A(a[49]), .B(b[49]), .Z(n21) );
  INV_X1 U124 ( .A(n84), .ZN(carry[4]) );
  AOI22_X1 U125 ( .A1(b[3]), .A2(a[3]), .B1(n31), .B2(c[3]), .ZN(n84) );
  XOR2_X1 U126 ( .A(a[3]), .B(b[3]), .Z(n31) );
  INV_X1 U127 ( .A(n85), .ZN(carry[49]) );
  AOI22_X1 U128 ( .A1(b[48]), .A2(a[48]), .B1(n22), .B2(c[48]), .ZN(n85) );
  XOR2_X1 U129 ( .A(a[48]), .B(b[48]), .Z(n22) );
  INV_X1 U130 ( .A(n86), .ZN(carry[48]) );
  AOI22_X1 U131 ( .A1(b[47]), .A2(a[47]), .B1(n23), .B2(c[47]), .ZN(n86) );
  XOR2_X1 U132 ( .A(a[47]), .B(b[47]), .Z(n23) );
  INV_X1 U133 ( .A(n87), .ZN(carry[47]) );
  AOI22_X1 U134 ( .A1(b[46]), .A2(a[46]), .B1(n24), .B2(c[46]), .ZN(n87) );
  XOR2_X1 U135 ( .A(a[46]), .B(b[46]), .Z(n24) );
  INV_X1 U136 ( .A(n88), .ZN(carry[46]) );
  AOI22_X1 U137 ( .A1(b[45]), .A2(a[45]), .B1(n25), .B2(c[45]), .ZN(n88) );
  XOR2_X1 U138 ( .A(a[45]), .B(b[45]), .Z(n25) );
  INV_X1 U139 ( .A(n89), .ZN(carry[45]) );
  AOI22_X1 U140 ( .A1(b[44]), .A2(a[44]), .B1(n26), .B2(c[44]), .ZN(n89) );
  XOR2_X1 U141 ( .A(a[44]), .B(b[44]), .Z(n26) );
  INV_X1 U142 ( .A(n90), .ZN(carry[44]) );
  AOI22_X1 U143 ( .A1(b[43]), .A2(a[43]), .B1(n27), .B2(c[43]), .ZN(n90) );
  XOR2_X1 U144 ( .A(a[43]), .B(b[43]), .Z(n27) );
  INV_X1 U145 ( .A(n91), .ZN(carry[43]) );
  AOI22_X1 U146 ( .A1(b[42]), .A2(a[42]), .B1(n28), .B2(c[42]), .ZN(n91) );
  XOR2_X1 U147 ( .A(a[42]), .B(b[42]), .Z(n28) );
  INV_X1 U148 ( .A(n92), .ZN(carry[42]) );
  AOI22_X1 U149 ( .A1(b[41]), .A2(a[41]), .B1(n29), .B2(c[41]), .ZN(n92) );
  XOR2_X1 U150 ( .A(a[41]), .B(b[41]), .Z(n29) );
  INV_X1 U151 ( .A(n93), .ZN(carry[41]) );
  AOI22_X1 U152 ( .A1(b[40]), .A2(a[40]), .B1(n30), .B2(c[40]), .ZN(n93) );
  XOR2_X1 U153 ( .A(a[40]), .B(b[40]), .Z(n30) );
  INV_X1 U154 ( .A(n94), .ZN(carry[40]) );
  AOI22_X1 U155 ( .A1(b[39]), .A2(a[39]), .B1(n32), .B2(c[39]), .ZN(n94) );
  XOR2_X1 U156 ( .A(a[39]), .B(b[39]), .Z(n32) );
  INV_X1 U157 ( .A(n95), .ZN(carry[3]) );
  AOI22_X1 U158 ( .A1(b[2]), .A2(a[2]), .B1(n42), .B2(c[2]), .ZN(n95) );
  XOR2_X1 U159 ( .A(a[2]), .B(b[2]), .Z(n42) );
  INV_X1 U160 ( .A(n96), .ZN(carry[39]) );
  AOI22_X1 U161 ( .A1(b[38]), .A2(a[38]), .B1(n33), .B2(c[38]), .ZN(n96) );
  XOR2_X1 U162 ( .A(a[38]), .B(b[38]), .Z(n33) );
  INV_X1 U163 ( .A(n97), .ZN(carry[38]) );
  AOI22_X1 U164 ( .A1(b[37]), .A2(a[37]), .B1(n34), .B2(c[37]), .ZN(n97) );
  XOR2_X1 U165 ( .A(a[37]), .B(b[37]), .Z(n34) );
  INV_X1 U166 ( .A(n98), .ZN(carry[37]) );
  AOI22_X1 U167 ( .A1(b[36]), .A2(a[36]), .B1(n35), .B2(c[36]), .ZN(n98) );
  XOR2_X1 U168 ( .A(a[36]), .B(b[36]), .Z(n35) );
  INV_X1 U169 ( .A(n99), .ZN(carry[36]) );
  AOI22_X1 U170 ( .A1(b[35]), .A2(a[35]), .B1(n36), .B2(c[35]), .ZN(n99) );
  XOR2_X1 U171 ( .A(a[35]), .B(b[35]), .Z(n36) );
  INV_X1 U172 ( .A(n100), .ZN(carry[35]) );
  AOI22_X1 U173 ( .A1(b[34]), .A2(a[34]), .B1(n37), .B2(c[34]), .ZN(n100) );
  XOR2_X1 U174 ( .A(a[34]), .B(b[34]), .Z(n37) );
  INV_X1 U175 ( .A(n101), .ZN(carry[34]) );
  AOI22_X1 U176 ( .A1(b[33]), .A2(a[33]), .B1(n38), .B2(c[33]), .ZN(n101) );
  XOR2_X1 U177 ( .A(a[33]), .B(b[33]), .Z(n38) );
  INV_X1 U178 ( .A(n102), .ZN(carry[33]) );
  AOI22_X1 U179 ( .A1(b[32]), .A2(a[32]), .B1(n39), .B2(c[32]), .ZN(n102) );
  XOR2_X1 U180 ( .A(a[32]), .B(b[32]), .Z(n39) );
  INV_X1 U181 ( .A(n103), .ZN(carry[32]) );
  AOI22_X1 U182 ( .A1(b[31]), .A2(a[31]), .B1(n40), .B2(c[31]), .ZN(n103) );
  XOR2_X1 U183 ( .A(a[31]), .B(b[31]), .Z(n40) );
  INV_X1 U184 ( .A(n104), .ZN(carry[31]) );
  AOI22_X1 U185 ( .A1(b[30]), .A2(a[30]), .B1(n41), .B2(c[30]), .ZN(n104) );
  XOR2_X1 U186 ( .A(a[30]), .B(b[30]), .Z(n41) );
  INV_X1 U187 ( .A(n105), .ZN(carry[30]) );
  AOI22_X1 U188 ( .A1(b[29]), .A2(a[29]), .B1(n43), .B2(c[29]), .ZN(n105) );
  XOR2_X1 U189 ( .A(a[29]), .B(b[29]), .Z(n43) );
  INV_X1 U190 ( .A(n106), .ZN(carry[2]) );
  AOI22_X1 U191 ( .A1(b[1]), .A2(a[1]), .B1(n53), .B2(c[1]), .ZN(n106) );
  XOR2_X1 U192 ( .A(a[1]), .B(b[1]), .Z(n53) );
  INV_X1 U193 ( .A(n107), .ZN(carry[29]) );
  AOI22_X1 U194 ( .A1(b[28]), .A2(a[28]), .B1(n44), .B2(c[28]), .ZN(n107) );
  XOR2_X1 U195 ( .A(a[28]), .B(b[28]), .Z(n44) );
  INV_X1 U196 ( .A(n108), .ZN(carry[28]) );
  AOI22_X1 U197 ( .A1(b[27]), .A2(a[27]), .B1(n45), .B2(c[27]), .ZN(n108) );
  XOR2_X1 U198 ( .A(a[27]), .B(b[27]), .Z(n45) );
  INV_X1 U199 ( .A(n109), .ZN(carry[27]) );
  AOI22_X1 U200 ( .A1(b[26]), .A2(a[26]), .B1(n46), .B2(c[26]), .ZN(n109) );
  XOR2_X1 U201 ( .A(a[26]), .B(b[26]), .Z(n46) );
  INV_X1 U202 ( .A(n110), .ZN(carry[26]) );
  AOI22_X1 U203 ( .A1(b[25]), .A2(a[25]), .B1(n47), .B2(c[25]), .ZN(n110) );
  XOR2_X1 U204 ( .A(a[25]), .B(b[25]), .Z(n47) );
  INV_X1 U205 ( .A(n111), .ZN(carry[25]) );
  AOI22_X1 U206 ( .A1(b[24]), .A2(a[24]), .B1(n48), .B2(c[24]), .ZN(n111) );
  XOR2_X1 U207 ( .A(a[24]), .B(b[24]), .Z(n48) );
  INV_X1 U208 ( .A(n112), .ZN(carry[24]) );
  AOI22_X1 U209 ( .A1(b[23]), .A2(a[23]), .B1(n49), .B2(c[23]), .ZN(n112) );
  XOR2_X1 U210 ( .A(a[23]), .B(b[23]), .Z(n49) );
  INV_X1 U211 ( .A(n113), .ZN(carry[23]) );
  AOI22_X1 U212 ( .A1(b[22]), .A2(a[22]), .B1(n50), .B2(c[22]), .ZN(n113) );
  XOR2_X1 U213 ( .A(a[22]), .B(b[22]), .Z(n50) );
  INV_X1 U214 ( .A(n114), .ZN(carry[22]) );
  AOI22_X1 U215 ( .A1(b[21]), .A2(a[21]), .B1(n51), .B2(c[21]), .ZN(n114) );
  XOR2_X1 U216 ( .A(a[21]), .B(b[21]), .Z(n51) );
  INV_X1 U217 ( .A(n115), .ZN(carry[21]) );
  AOI22_X1 U218 ( .A1(b[20]), .A2(a[20]), .B1(n52), .B2(c[20]), .ZN(n115) );
  XOR2_X1 U219 ( .A(a[20]), .B(b[20]), .Z(n52) );
  INV_X1 U220 ( .A(n116), .ZN(carry[20]) );
  AOI22_X1 U221 ( .A1(b[19]), .A2(a[19]), .B1(n54), .B2(c[19]), .ZN(n116) );
  XOR2_X1 U222 ( .A(a[19]), .B(b[19]), .Z(n54) );
  INV_X1 U223 ( .A(n117), .ZN(carry[1]) );
  AOI22_X1 U224 ( .A1(b[0]), .A2(a[0]), .B1(n64), .B2(c[0]), .ZN(n117) );
  XOR2_X1 U225 ( .A(a[0]), .B(b[0]), .Z(n64) );
  INV_X1 U226 ( .A(n118), .ZN(carry[19]) );
  AOI22_X1 U227 ( .A1(b[18]), .A2(a[18]), .B1(n55), .B2(c[18]), .ZN(n118) );
  XOR2_X1 U228 ( .A(a[18]), .B(b[18]), .Z(n55) );
  INV_X1 U229 ( .A(n119), .ZN(carry[18]) );
  AOI22_X1 U230 ( .A1(b[17]), .A2(a[17]), .B1(n56), .B2(c[17]), .ZN(n119) );
  XOR2_X1 U231 ( .A(a[17]), .B(b[17]), .Z(n56) );
  INV_X1 U232 ( .A(n120), .ZN(carry[17]) );
  AOI22_X1 U233 ( .A1(b[16]), .A2(a[16]), .B1(n57), .B2(c[16]), .ZN(n120) );
  XOR2_X1 U234 ( .A(a[16]), .B(b[16]), .Z(n57) );
  INV_X1 U235 ( .A(n121), .ZN(carry[16]) );
  AOI22_X1 U236 ( .A1(b[15]), .A2(a[15]), .B1(n58), .B2(c[15]), .ZN(n121) );
  XOR2_X1 U237 ( .A(a[15]), .B(b[15]), .Z(n58) );
  INV_X1 U238 ( .A(n122), .ZN(carry[15]) );
  AOI22_X1 U239 ( .A1(b[14]), .A2(a[14]), .B1(n59), .B2(c[14]), .ZN(n122) );
  XOR2_X1 U240 ( .A(a[14]), .B(b[14]), .Z(n59) );
  INV_X1 U241 ( .A(n123), .ZN(carry[14]) );
  AOI22_X1 U242 ( .A1(b[13]), .A2(a[13]), .B1(n60), .B2(c[13]), .ZN(n123) );
  XOR2_X1 U243 ( .A(a[13]), .B(b[13]), .Z(n60) );
  INV_X1 U244 ( .A(n124), .ZN(carry[13]) );
  AOI22_X1 U245 ( .A1(b[12]), .A2(a[12]), .B1(n61), .B2(c[12]), .ZN(n124) );
  XOR2_X1 U246 ( .A(a[12]), .B(b[12]), .Z(n61) );
  INV_X1 U247 ( .A(n125), .ZN(carry[12]) );
  AOI22_X1 U248 ( .A1(b[11]), .A2(a[11]), .B1(n62), .B2(c[11]), .ZN(n125) );
  XOR2_X1 U249 ( .A(a[11]), .B(b[11]), .Z(n62) );
  INV_X1 U250 ( .A(n126), .ZN(carry[11]) );
  AOI22_X1 U251 ( .A1(b[10]), .A2(a[10]), .B1(n63), .B2(c[10]), .ZN(n126) );
  XOR2_X1 U252 ( .A(a[10]), .B(b[10]), .Z(n63) );
  INV_X1 U253 ( .A(n127), .ZN(carry[10]) );
  AOI22_X1 U254 ( .A1(b[9]), .A2(a[9]), .B1(n1), .B2(c[9]), .ZN(n127) );
  XOR2_X1 U255 ( .A(a[9]), .B(b[9]), .Z(n1) );
endmodule


module TM ( a, b, result );
  input [31:0] a;
  input [31:0] b;
  output [63:0] result;
  wire   shiftedA_7__37_, shiftedA_7__36_, shiftedA_7__35_, shiftedA_7__34_,
         shiftedA_7__33_, shiftedA_7__32_, shiftedA_7__31_, shiftedA_7__30_,
         shiftedA_7__29_, shiftedA_7__28_, shiftedA_7__27_, shiftedA_7__26_,
         shiftedA_7__25_, shiftedA_7__24_, shiftedA_7__23_, shiftedA_7__22_,
         shiftedA_7__21_, shiftedA_7__20_, shiftedA_7__19_, shiftedA_7__18_,
         shiftedA_7__17_, shiftedA_7__16_, shiftedA_7__15_, shiftedA_7__14_,
         shiftedA_7__13_, shiftedA_7__12_, shiftedA_7__11_, shiftedA_7__10_,
         shiftedA_7__9_, shiftedA_7__8_, shiftedA_7__7_, shiftedA_6__36_,
         shiftedA_6__35_, shiftedA_6__34_, shiftedA_6__33_, shiftedA_6__32_,
         shiftedA_6__31_, shiftedA_6__30_, shiftedA_6__29_, shiftedA_6__28_,
         shiftedA_6__27_, shiftedA_6__26_, shiftedA_6__25_, shiftedA_6__24_,
         shiftedA_6__23_, shiftedA_6__22_, shiftedA_6__21_, shiftedA_6__20_,
         shiftedA_6__19_, shiftedA_6__18_, shiftedA_6__17_, shiftedA_6__16_,
         shiftedA_6__15_, shiftedA_6__14_, shiftedA_6__13_, shiftedA_6__12_,
         shiftedA_6__11_, shiftedA_6__10_, shiftedA_6__9_, shiftedA_6__8_,
         shiftedA_6__7_, shiftedA_6__6_, shiftedA_5__35_, shiftedA_5__34_,
         shiftedA_5__33_, shiftedA_5__32_, shiftedA_5__31_, shiftedA_5__30_,
         shiftedA_5__29_, shiftedA_5__28_, shiftedA_5__27_, shiftedA_5__26_,
         shiftedA_5__25_, shiftedA_5__24_, shiftedA_5__23_, shiftedA_5__22_,
         shiftedA_5__21_, shiftedA_5__20_, shiftedA_5__19_, shiftedA_5__18_,
         shiftedA_5__17_, shiftedA_5__16_, shiftedA_5__15_, shiftedA_5__14_,
         shiftedA_5__13_, shiftedA_5__12_, shiftedA_5__11_, shiftedA_5__10_,
         shiftedA_5__9_, shiftedA_5__8_, shiftedA_5__7_, shiftedA_5__6_,
         shiftedA_5__5_, shiftedA_4__34_, shiftedA_4__33_, shiftedA_4__32_,
         shiftedA_4__31_, shiftedA_4__30_, shiftedA_4__29_, shiftedA_4__28_,
         shiftedA_4__27_, shiftedA_4__26_, shiftedA_4__25_, shiftedA_4__24_,
         shiftedA_4__23_, shiftedA_4__22_, shiftedA_4__21_, shiftedA_4__20_,
         shiftedA_4__19_, shiftedA_4__18_, shiftedA_4__17_, shiftedA_4__16_,
         shiftedA_4__15_, shiftedA_4__14_, shiftedA_4__13_, shiftedA_4__12_,
         shiftedA_4__11_, shiftedA_4__10_, shiftedA_4__9_, shiftedA_4__8_,
         shiftedA_4__7_, shiftedA_4__6_, shiftedA_4__5_, shiftedA_4__4_,
         shiftedA_3__33_, shiftedA_3__32_, shiftedA_3__31_, shiftedA_3__30_,
         shiftedA_3__29_, shiftedA_3__28_, shiftedA_3__27_, shiftedA_3__26_,
         shiftedA_3__25_, shiftedA_3__24_, shiftedA_3__23_, shiftedA_3__22_,
         shiftedA_3__21_, shiftedA_3__20_, shiftedA_3__19_, shiftedA_3__18_,
         shiftedA_3__17_, shiftedA_3__16_, shiftedA_3__15_, shiftedA_3__14_,
         shiftedA_3__13_, shiftedA_3__12_, shiftedA_3__11_, shiftedA_3__10_,
         shiftedA_3__9_, shiftedA_3__8_, shiftedA_3__7_, shiftedA_3__6_,
         shiftedA_3__5_, shiftedA_3__4_, shiftedA_3__3_, shiftedA_2__32_,
         shiftedA_2__31_, shiftedA_2__30_, shiftedA_2__29_, shiftedA_2__28_,
         shiftedA_2__27_, shiftedA_2__26_, shiftedA_2__25_, shiftedA_2__24_,
         shiftedA_2__23_, shiftedA_2__22_, shiftedA_2__21_, shiftedA_2__20_,
         shiftedA_2__19_, shiftedA_2__18_, shiftedA_2__17_, shiftedA_2__16_,
         shiftedA_2__15_, shiftedA_2__14_, shiftedA_2__13_, shiftedA_2__12_,
         shiftedA_2__11_, shiftedA_2__10_, shiftedA_2__9_, shiftedA_2__8_,
         shiftedA_2__7_, shiftedA_2__6_, shiftedA_2__5_, shiftedA_2__4_,
         shiftedA_2__3_, shiftedA_2__2_, shiftedA_1__31_, shiftedA_1__30_,
         shiftedA_1__29_, shiftedA_1__28_, shiftedA_1__27_, shiftedA_1__26_,
         shiftedA_1__25_, shiftedA_1__24_, shiftedA_1__23_, shiftedA_1__22_,
         shiftedA_1__21_, shiftedA_1__20_, shiftedA_1__19_, shiftedA_1__18_,
         shiftedA_1__17_, shiftedA_1__16_, shiftedA_1__15_, shiftedA_1__14_,
         shiftedA_1__13_, shiftedA_1__12_, shiftedA_1__11_, shiftedA_1__10_,
         shiftedA_1__9_, shiftedA_1__8_, shiftedA_1__7_, shiftedA_1__6_,
         shiftedA_1__5_, shiftedA_1__4_, shiftedA_1__3_, shiftedA_1__2_,
         shiftedA_1__1_, shiftedA_0__30_, shiftedA_0__29_, shiftedA_0__28_,
         shiftedA_0__27_, shiftedA_0__26_, shiftedA_0__25_, shiftedA_0__24_,
         shiftedA_0__23_, shiftedA_0__22_, shiftedA_0__21_, shiftedA_0__20_,
         shiftedA_0__19_, shiftedA_0__18_, shiftedA_0__17_, shiftedA_0__16_,
         shiftedA_0__15_, shiftedA_0__14_, shiftedA_0__13_, shiftedA_0__12_,
         shiftedA_0__11_, shiftedA_0__10_, shiftedA_0__9_, shiftedA_0__8_,
         shiftedA_0__7_, shiftedA_0__6_, shiftedA_0__5_, shiftedA_0__4_,
         shiftedA_0__3_, shiftedA_0__2_, shiftedA_0__1_, shiftedA_0__0_,
         shiftedA_45__63_, shiftedA_44__63_, shiftedA_43__63_,
         shiftedA_42__63_, shiftedA_41__63_, shiftedA_40__63_,
         shiftedA_39__63_, shiftedA_38__63_, shiftedA_37__63_,
         shiftedA_36__63_, shiftedA_35__63_, shiftedA_34__63_,
         shiftedA_33__63_, shiftedA_32__63_, shiftedA_30__63_,
         shiftedA_30__60_, shiftedA_30__59_, shiftedA_30__58_,
         shiftedA_30__57_, shiftedA_30__56_, shiftedA_30__55_,
         shiftedA_30__54_, shiftedA_30__53_, shiftedA_30__52_,
         shiftedA_30__51_, shiftedA_30__50_, shiftedA_30__49_,
         shiftedA_30__48_, shiftedA_30__47_, shiftedA_30__46_,
         shiftedA_30__45_, shiftedA_30__44_, shiftedA_30__43_,
         shiftedA_30__42_, shiftedA_30__41_, shiftedA_30__40_,
         shiftedA_30__39_, shiftedA_30__38_, shiftedA_30__37_,
         shiftedA_30__36_, shiftedA_30__35_, shiftedA_30__34_,
         shiftedA_30__33_, shiftedA_30__32_, shiftedA_30__31_,
         shiftedA_30__30_, shiftedA_29__63_, shiftedA_29__59_,
         shiftedA_29__58_, shiftedA_29__57_, shiftedA_29__56_,
         shiftedA_29__55_, shiftedA_29__54_, shiftedA_29__53_,
         shiftedA_29__52_, shiftedA_29__51_, shiftedA_29__50_,
         shiftedA_29__49_, shiftedA_29__48_, shiftedA_29__47_,
         shiftedA_29__46_, shiftedA_29__45_, shiftedA_29__44_,
         shiftedA_29__43_, shiftedA_29__42_, shiftedA_29__41_,
         shiftedA_29__40_, shiftedA_29__39_, shiftedA_29__38_,
         shiftedA_29__37_, shiftedA_29__36_, shiftedA_29__35_,
         shiftedA_29__34_, shiftedA_29__33_, shiftedA_29__32_,
         shiftedA_29__31_, shiftedA_29__30_, shiftedA_29__29_,
         shiftedA_28__63_, shiftedA_28__58_, shiftedA_28__57_,
         shiftedA_28__56_, shiftedA_28__55_, shiftedA_28__54_,
         shiftedA_28__53_, shiftedA_28__52_, shiftedA_28__51_,
         shiftedA_28__50_, shiftedA_28__49_, shiftedA_28__48_,
         shiftedA_28__47_, shiftedA_28__46_, shiftedA_28__45_,
         shiftedA_28__44_, shiftedA_28__43_, shiftedA_28__42_,
         shiftedA_28__41_, shiftedA_28__40_, shiftedA_28__39_,
         shiftedA_28__38_, shiftedA_28__37_, shiftedA_28__36_,
         shiftedA_28__35_, shiftedA_28__34_, shiftedA_28__33_,
         shiftedA_28__32_, shiftedA_28__31_, shiftedA_28__30_,
         shiftedA_28__29_, shiftedA_28__28_, shiftedA_27__63_,
         shiftedA_27__57_, shiftedA_27__56_, shiftedA_27__55_,
         shiftedA_27__54_, shiftedA_27__53_, shiftedA_27__52_,
         shiftedA_27__51_, shiftedA_27__50_, shiftedA_27__49_,
         shiftedA_27__48_, shiftedA_27__47_, shiftedA_27__46_,
         shiftedA_27__45_, shiftedA_27__44_, shiftedA_27__43_,
         shiftedA_27__42_, shiftedA_27__41_, shiftedA_27__40_,
         shiftedA_27__39_, shiftedA_27__38_, shiftedA_27__37_,
         shiftedA_27__36_, shiftedA_27__35_, shiftedA_27__34_,
         shiftedA_27__33_, shiftedA_27__32_, shiftedA_27__31_,
         shiftedA_27__30_, shiftedA_27__29_, shiftedA_27__28_,
         shiftedA_27__27_, shiftedA_26__63_, shiftedA_26__56_,
         shiftedA_26__55_, shiftedA_26__54_, shiftedA_26__53_,
         shiftedA_26__52_, shiftedA_26__51_, shiftedA_26__50_,
         shiftedA_26__49_, shiftedA_26__48_, shiftedA_26__47_,
         shiftedA_26__46_, shiftedA_26__45_, shiftedA_26__44_,
         shiftedA_26__43_, shiftedA_26__42_, shiftedA_26__41_,
         shiftedA_26__40_, shiftedA_26__39_, shiftedA_26__38_,
         shiftedA_26__37_, shiftedA_26__36_, shiftedA_26__35_,
         shiftedA_26__34_, shiftedA_26__33_, shiftedA_26__32_,
         shiftedA_26__31_, shiftedA_26__30_, shiftedA_26__29_,
         shiftedA_26__28_, shiftedA_26__27_, shiftedA_26__26_,
         shiftedA_25__63_, shiftedA_25__55_, shiftedA_25__54_,
         shiftedA_25__53_, shiftedA_25__52_, shiftedA_25__51_,
         shiftedA_25__50_, shiftedA_25__49_, shiftedA_25__48_,
         shiftedA_25__47_, shiftedA_25__46_, shiftedA_25__45_,
         shiftedA_25__44_, shiftedA_25__43_, shiftedA_25__42_,
         shiftedA_25__41_, shiftedA_25__40_, shiftedA_25__39_,
         shiftedA_25__38_, shiftedA_25__37_, shiftedA_25__36_,
         shiftedA_25__35_, shiftedA_25__34_, shiftedA_25__33_,
         shiftedA_25__32_, shiftedA_25__31_, shiftedA_25__30_,
         shiftedA_25__29_, shiftedA_25__28_, shiftedA_25__27_,
         shiftedA_25__26_, shiftedA_25__25_, shiftedA_24__63_,
         shiftedA_24__54_, shiftedA_24__53_, shiftedA_24__52_,
         shiftedA_24__51_, shiftedA_24__50_, shiftedA_24__49_,
         shiftedA_24__48_, shiftedA_24__47_, shiftedA_24__46_,
         shiftedA_24__45_, shiftedA_24__44_, shiftedA_24__43_,
         shiftedA_24__42_, shiftedA_24__41_, shiftedA_24__40_,
         shiftedA_24__39_, shiftedA_24__38_, shiftedA_24__37_,
         shiftedA_24__36_, shiftedA_24__35_, shiftedA_24__34_,
         shiftedA_24__33_, shiftedA_24__32_, shiftedA_24__31_,
         shiftedA_24__30_, shiftedA_24__29_, shiftedA_24__28_,
         shiftedA_24__27_, shiftedA_24__26_, shiftedA_24__25_,
         shiftedA_24__24_, shiftedA_23__63_, shiftedA_23__53_,
         shiftedA_23__52_, shiftedA_23__51_, shiftedA_23__50_,
         shiftedA_23__49_, shiftedA_23__48_, shiftedA_23__47_,
         shiftedA_23__46_, shiftedA_23__45_, shiftedA_23__44_,
         shiftedA_23__43_, shiftedA_23__42_, shiftedA_23__41_,
         shiftedA_23__40_, shiftedA_23__39_, shiftedA_23__38_,
         shiftedA_23__37_, shiftedA_23__36_, shiftedA_23__35_,
         shiftedA_23__34_, shiftedA_23__33_, shiftedA_23__32_,
         shiftedA_23__31_, shiftedA_23__30_, shiftedA_23__29_,
         shiftedA_23__28_, shiftedA_23__27_, shiftedA_23__26_,
         shiftedA_23__25_, shiftedA_23__24_, shiftedA_23__23_,
         shiftedA_22__63_, shiftedA_22__52_, shiftedA_22__51_,
         shiftedA_22__50_, shiftedA_22__49_, shiftedA_22__48_,
         shiftedA_22__47_, shiftedA_22__46_, shiftedA_22__45_,
         shiftedA_22__44_, shiftedA_22__43_, shiftedA_22__42_,
         shiftedA_22__41_, shiftedA_22__40_, shiftedA_22__39_,
         shiftedA_22__38_, shiftedA_22__37_, shiftedA_22__36_,
         shiftedA_22__35_, shiftedA_22__34_, shiftedA_22__33_,
         shiftedA_22__32_, shiftedA_22__31_, shiftedA_22__30_,
         shiftedA_22__29_, shiftedA_22__28_, shiftedA_22__27_,
         shiftedA_22__26_, shiftedA_22__25_, shiftedA_22__24_,
         shiftedA_22__23_, shiftedA_22__22_, shiftedA_21__63_,
         shiftedA_21__51_, shiftedA_21__50_, shiftedA_21__49_,
         shiftedA_21__48_, shiftedA_21__47_, shiftedA_21__46_,
         shiftedA_21__45_, shiftedA_21__44_, shiftedA_21__43_,
         shiftedA_21__42_, shiftedA_21__41_, shiftedA_21__40_,
         shiftedA_21__39_, shiftedA_21__38_, shiftedA_21__37_,
         shiftedA_21__36_, shiftedA_21__35_, shiftedA_21__34_,
         shiftedA_21__33_, shiftedA_21__32_, shiftedA_21__31_,
         shiftedA_21__30_, shiftedA_21__29_, shiftedA_21__28_,
         shiftedA_21__27_, shiftedA_21__26_, shiftedA_21__25_,
         shiftedA_21__24_, shiftedA_21__23_, shiftedA_21__22_,
         shiftedA_21__21_, shiftedA_20__63_, shiftedA_20__50_,
         shiftedA_20__49_, shiftedA_20__48_, shiftedA_20__47_,
         shiftedA_20__46_, shiftedA_20__45_, shiftedA_20__44_,
         shiftedA_20__43_, shiftedA_20__42_, shiftedA_20__41_,
         shiftedA_20__40_, shiftedA_20__39_, shiftedA_20__38_,
         shiftedA_20__37_, shiftedA_20__36_, shiftedA_20__35_,
         shiftedA_20__34_, shiftedA_20__33_, shiftedA_20__32_,
         shiftedA_20__31_, shiftedA_20__30_, shiftedA_20__29_,
         shiftedA_20__28_, shiftedA_20__27_, shiftedA_20__26_,
         shiftedA_20__25_, shiftedA_20__24_, shiftedA_20__23_,
         shiftedA_20__22_, shiftedA_20__21_, shiftedA_20__20_,
         shiftedA_19__63_, shiftedA_19__49_, shiftedA_19__48_,
         shiftedA_19__47_, shiftedA_19__46_, shiftedA_19__45_,
         shiftedA_19__44_, shiftedA_19__43_, shiftedA_19__42_,
         shiftedA_19__41_, shiftedA_19__40_, shiftedA_19__39_,
         shiftedA_19__38_, shiftedA_19__37_, shiftedA_19__36_,
         shiftedA_19__35_, shiftedA_19__34_, shiftedA_19__33_,
         shiftedA_19__32_, shiftedA_19__31_, shiftedA_19__30_,
         shiftedA_19__29_, shiftedA_19__28_, shiftedA_19__27_,
         shiftedA_19__26_, shiftedA_19__25_, shiftedA_19__24_,
         shiftedA_19__23_, shiftedA_19__22_, shiftedA_19__21_,
         shiftedA_19__20_, shiftedA_19__19_, shiftedA_18__63_,
         shiftedA_18__48_, shiftedA_18__47_, shiftedA_18__46_,
         shiftedA_18__45_, shiftedA_18__44_, shiftedA_18__43_,
         shiftedA_18__42_, shiftedA_18__41_, shiftedA_18__40_,
         shiftedA_18__39_, shiftedA_18__38_, shiftedA_18__37_,
         shiftedA_18__36_, shiftedA_18__35_, shiftedA_18__34_,
         shiftedA_18__33_, shiftedA_18__32_, shiftedA_18__31_,
         shiftedA_18__30_, shiftedA_18__29_, shiftedA_18__28_,
         shiftedA_18__27_, shiftedA_18__26_, shiftedA_18__25_,
         shiftedA_18__24_, shiftedA_18__23_, shiftedA_18__22_,
         shiftedA_18__21_, shiftedA_18__20_, shiftedA_18__19_,
         shiftedA_18__18_, shiftedA_17__47_, shiftedA_17__46_,
         shiftedA_17__45_, shiftedA_17__44_, shiftedA_17__43_,
         shiftedA_17__42_, shiftedA_17__41_, shiftedA_17__40_,
         shiftedA_17__39_, shiftedA_17__38_, shiftedA_17__37_,
         shiftedA_17__36_, shiftedA_17__35_, shiftedA_17__34_,
         shiftedA_17__33_, shiftedA_17__32_, shiftedA_17__31_,
         shiftedA_17__30_, shiftedA_17__29_, shiftedA_17__28_,
         shiftedA_17__27_, shiftedA_17__26_, shiftedA_17__25_,
         shiftedA_17__24_, shiftedA_17__23_, shiftedA_17__22_,
         shiftedA_17__21_, shiftedA_17__20_, shiftedA_17__19_,
         shiftedA_17__18_, shiftedA_17__17_, shiftedA_16__46_,
         shiftedA_16__45_, shiftedA_16__44_, shiftedA_16__43_,
         shiftedA_16__42_, shiftedA_16__41_, shiftedA_16__40_,
         shiftedA_16__39_, shiftedA_16__38_, shiftedA_16__37_,
         shiftedA_16__36_, shiftedA_16__35_, shiftedA_16__34_,
         shiftedA_16__33_, shiftedA_16__32_, shiftedA_16__31_,
         shiftedA_16__30_, shiftedA_16__29_, shiftedA_16__28_,
         shiftedA_16__27_, shiftedA_16__26_, shiftedA_16__25_,
         shiftedA_16__24_, shiftedA_16__23_, shiftedA_16__22_,
         shiftedA_16__21_, shiftedA_16__20_, shiftedA_16__19_,
         shiftedA_16__18_, shiftedA_16__17_, shiftedA_16__16_,
         shiftedA_15__45_, shiftedA_15__44_, shiftedA_15__43_,
         shiftedA_15__42_, shiftedA_15__41_, shiftedA_15__40_,
         shiftedA_15__39_, shiftedA_15__38_, shiftedA_15__37_,
         shiftedA_15__36_, shiftedA_15__35_, shiftedA_15__34_,
         shiftedA_15__33_, shiftedA_15__32_, shiftedA_15__31_,
         shiftedA_15__30_, shiftedA_15__29_, shiftedA_15__28_,
         shiftedA_15__27_, shiftedA_15__26_, shiftedA_15__25_,
         shiftedA_15__24_, shiftedA_15__23_, shiftedA_15__22_,
         shiftedA_15__21_, shiftedA_15__20_, shiftedA_15__19_,
         shiftedA_15__18_, shiftedA_15__17_, shiftedA_15__16_,
         shiftedA_15__15_, shiftedA_14__44_, shiftedA_14__43_,
         shiftedA_14__42_, shiftedA_14__41_, shiftedA_14__40_,
         shiftedA_14__39_, shiftedA_14__38_, shiftedA_14__37_,
         shiftedA_14__36_, shiftedA_14__35_, shiftedA_14__34_,
         shiftedA_14__33_, shiftedA_14__32_, shiftedA_14__31_,
         shiftedA_14__30_, shiftedA_14__29_, shiftedA_14__28_,
         shiftedA_14__27_, shiftedA_14__26_, shiftedA_14__25_,
         shiftedA_14__24_, shiftedA_14__23_, shiftedA_14__22_,
         shiftedA_14__21_, shiftedA_14__20_, shiftedA_14__19_,
         shiftedA_14__18_, shiftedA_14__17_, shiftedA_14__16_,
         shiftedA_14__15_, shiftedA_14__14_, shiftedA_13__43_,
         shiftedA_13__42_, shiftedA_13__41_, shiftedA_13__40_,
         shiftedA_13__39_, shiftedA_13__38_, shiftedA_13__37_,
         shiftedA_13__36_, shiftedA_13__35_, shiftedA_13__34_,
         shiftedA_13__33_, shiftedA_13__32_, shiftedA_13__31_,
         shiftedA_13__30_, shiftedA_13__29_, shiftedA_13__28_,
         shiftedA_13__27_, shiftedA_13__26_, shiftedA_13__25_,
         shiftedA_13__24_, shiftedA_13__23_, shiftedA_13__22_,
         shiftedA_13__21_, shiftedA_13__20_, shiftedA_13__19_,
         shiftedA_13__18_, shiftedA_13__17_, shiftedA_13__16_,
         shiftedA_13__15_, shiftedA_13__14_, shiftedA_13__13_,
         shiftedA_12__42_, shiftedA_12__41_, shiftedA_12__40_,
         shiftedA_12__39_, shiftedA_12__38_, shiftedA_12__37_,
         shiftedA_12__36_, shiftedA_12__35_, shiftedA_12__34_,
         shiftedA_12__33_, shiftedA_12__32_, shiftedA_12__31_,
         shiftedA_12__30_, shiftedA_12__29_, shiftedA_12__28_,
         shiftedA_12__27_, shiftedA_12__26_, shiftedA_12__25_,
         shiftedA_12__24_, shiftedA_12__23_, shiftedA_12__22_,
         shiftedA_12__21_, shiftedA_12__20_, shiftedA_12__19_,
         shiftedA_12__18_, shiftedA_12__17_, shiftedA_12__16_,
         shiftedA_12__15_, shiftedA_12__14_, shiftedA_12__13_,
         shiftedA_12__12_, shiftedA_11__41_, shiftedA_11__40_,
         shiftedA_11__39_, shiftedA_11__38_, shiftedA_11__37_,
         shiftedA_11__36_, shiftedA_11__35_, shiftedA_11__34_,
         shiftedA_11__33_, shiftedA_11__32_, shiftedA_11__31_,
         shiftedA_11__30_, shiftedA_11__29_, shiftedA_11__28_,
         shiftedA_11__27_, shiftedA_11__26_, shiftedA_11__25_,
         shiftedA_11__24_, shiftedA_11__23_, shiftedA_11__22_,
         shiftedA_11__21_, shiftedA_11__20_, shiftedA_11__19_,
         shiftedA_11__18_, shiftedA_11__17_, shiftedA_11__16_,
         shiftedA_11__15_, shiftedA_11__14_, shiftedA_11__13_,
         shiftedA_11__12_, shiftedA_11__11_, shiftedA_10__40_,
         shiftedA_10__39_, shiftedA_10__38_, shiftedA_10__37_,
         shiftedA_10__36_, shiftedA_10__35_, shiftedA_10__34_,
         shiftedA_10__33_, shiftedA_10__32_, shiftedA_10__31_,
         shiftedA_10__30_, shiftedA_10__29_, shiftedA_10__28_,
         shiftedA_10__27_, shiftedA_10__26_, shiftedA_10__25_,
         shiftedA_10__24_, shiftedA_10__23_, shiftedA_10__22_,
         shiftedA_10__21_, shiftedA_10__20_, shiftedA_10__19_,
         shiftedA_10__18_, shiftedA_10__17_, shiftedA_10__16_,
         shiftedA_10__15_, shiftedA_10__14_, shiftedA_10__13_,
         shiftedA_10__12_, shiftedA_10__11_, shiftedA_10__10_, shiftedA_9__39_,
         shiftedA_9__38_, shiftedA_9__37_, shiftedA_9__36_, shiftedA_9__35_,
         shiftedA_9__34_, shiftedA_9__33_, shiftedA_9__32_, shiftedA_9__31_,
         shiftedA_9__30_, shiftedA_9__29_, shiftedA_9__28_, shiftedA_9__27_,
         shiftedA_9__26_, shiftedA_9__25_, shiftedA_9__24_, shiftedA_9__23_,
         shiftedA_9__22_, shiftedA_9__21_, shiftedA_9__20_, shiftedA_9__19_,
         shiftedA_9__18_, shiftedA_9__17_, shiftedA_9__16_, shiftedA_9__15_,
         shiftedA_9__14_, shiftedA_9__13_, shiftedA_9__12_, shiftedA_9__11_,
         shiftedA_9__10_, shiftedA_9__9_, shiftedA_8__38_, shiftedA_8__37_,
         shiftedA_8__36_, shiftedA_8__35_, shiftedA_8__34_, shiftedA_8__33_,
         shiftedA_8__32_, shiftedA_8__31_, shiftedA_8__30_, shiftedA_8__29_,
         shiftedA_8__28_, shiftedA_8__27_, shiftedA_8__26_, shiftedA_8__25_,
         shiftedA_8__24_, shiftedA_8__23_, shiftedA_8__22_, shiftedA_8__21_,
         shiftedA_8__20_, shiftedA_8__19_, shiftedA_8__18_, shiftedA_8__17_,
         shiftedA_8__16_, shiftedA_8__15_, shiftedA_8__14_, shiftedA_8__13_,
         shiftedA_8__12_, shiftedA_8__11_, shiftedA_8__10_, shiftedA_8__9_,
         shiftedA_8__8_, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199;
  wire   [1343:0] adderResult_level1;
  wire   [1343:0] carry_level1;
  wire   [895:0] adderResult_level2;
  wire   [895:0] carry_level2;
  wire   [575:0] adderResult_level3;
  wire   [575:0] carry_level3;
  wire   [383:0] adderResult_level4;
  wire   [383:0] carry_level4;
  wire   [255:0] adderResult_level5;
  wire   [255:0] carry_level5;
  wire   [191:0] adderResult_level6;
  wire   [191:0] carry_level6;
  wire   [127:0] adderResult_level7;
  wire   [127:0] carry_level7;
  wire   [63:0] adderResult_level8;
  wire   [63:0] carry_level8;
  wire   [63:0] adderResult_level9;
  wire   [63:0] carry_level9;
  wire   [63:0] adderResult_level10;
  wire   [63:0] carry_level10;

  BWAdder_0 level1_0__adder ( .a({n134, n134, n134, n134, n134, n134, n134, 
        n134, n134, n134, n134, n134, n134, n134, n134, n134, n134, n134, n134, 
        n134, n134, n134, n134, n134, n134, n134, n134, n134, n134, n134, n134, 
        n134, n134, shiftedA_0__30_, shiftedA_0__29_, shiftedA_0__28_, 
        shiftedA_0__27_, shiftedA_0__26_, shiftedA_0__25_, shiftedA_0__24_, 
        shiftedA_0__23_, shiftedA_0__22_, shiftedA_0__21_, shiftedA_0__20_, 
        shiftedA_0__19_, shiftedA_0__18_, shiftedA_0__17_, shiftedA_0__16_, 
        shiftedA_0__15_, shiftedA_0__14_, shiftedA_0__13_, shiftedA_0__12_, 
        shiftedA_0__11_, shiftedA_0__10_, shiftedA_0__9_, shiftedA_0__8_, 
        shiftedA_0__7_, shiftedA_0__6_, shiftedA_0__5_, shiftedA_0__4_, 
        shiftedA_0__3_, shiftedA_0__2_, shiftedA_0__1_, shiftedA_0__0_}), .b({
        n131, n131, n131, n131, n131, n131, n131, n131, n131, n131, n131, n131, 
        n131, n131, n131, n131, n131, n131, n131, n131, n131, n131, n131, n131, 
        n131, n131, n131, n131, n131, n131, n131, n131, shiftedA_1__31_, 
        shiftedA_1__30_, shiftedA_1__29_, shiftedA_1__28_, shiftedA_1__27_, 
        shiftedA_1__26_, shiftedA_1__25_, shiftedA_1__24_, shiftedA_1__23_, 
        shiftedA_1__22_, shiftedA_1__21_, shiftedA_1__20_, shiftedA_1__19_, 
        shiftedA_1__18_, shiftedA_1__17_, shiftedA_1__16_, shiftedA_1__15_, 
        shiftedA_1__14_, shiftedA_1__13_, shiftedA_1__12_, shiftedA_1__11_, 
        shiftedA_1__10_, shiftedA_1__9_, shiftedA_1__8_, shiftedA_1__7_, 
        shiftedA_1__6_, shiftedA_1__5_, shiftedA_1__4_, shiftedA_1__3_, 
        shiftedA_1__2_, shiftedA_1__1_, 1'b0}), .c({n130, n130, n130, n130, 
        n130, n130, n130, n130, n130, n130, n130, n130, n130, n130, n130, n130, 
        n130, n130, n130, n130, n130, n130, n130, n130, n130, n130, n130, n130, 
        n130, n130, n130, shiftedA_2__32_, shiftedA_2__31_, shiftedA_2__30_, 
        shiftedA_2__29_, shiftedA_2__28_, shiftedA_2__27_, shiftedA_2__26_, 
        shiftedA_2__25_, shiftedA_2__24_, shiftedA_2__23_, shiftedA_2__22_, 
        shiftedA_2__21_, shiftedA_2__20_, shiftedA_2__19_, shiftedA_2__18_, 
        shiftedA_2__17_, shiftedA_2__16_, shiftedA_2__15_, shiftedA_2__14_, 
        shiftedA_2__13_, shiftedA_2__12_, shiftedA_2__11_, shiftedA_2__10_, 
        shiftedA_2__9_, shiftedA_2__8_, shiftedA_2__7_, shiftedA_2__6_, 
        shiftedA_2__5_, shiftedA_2__4_, shiftedA_2__3_, shiftedA_2__2_, 1'b0, 
        1'b0}), .result(adderResult_level1[63:0]), .carry(carry_level1[63:0])
         );
  BWAdder_61 level1_1__adder ( .a({n128, n128, n128, n128, n128, n128, n128, 
        n128, n128, n128, n128, n128, n128, n128, n128, n128, n128, n128, n128, 
        n128, n128, n128, n128, n128, n128, n128, n128, n128, n128, n128, 
        shiftedA_3__33_, shiftedA_3__32_, shiftedA_3__31_, shiftedA_3__30_, 
        shiftedA_3__29_, shiftedA_3__28_, shiftedA_3__27_, shiftedA_3__26_, 
        shiftedA_3__25_, shiftedA_3__24_, shiftedA_3__23_, shiftedA_3__22_, 
        shiftedA_3__21_, shiftedA_3__20_, shiftedA_3__19_, shiftedA_3__18_, 
        shiftedA_3__17_, shiftedA_3__16_, shiftedA_3__15_, shiftedA_3__14_, 
        shiftedA_3__13_, shiftedA_3__12_, shiftedA_3__11_, shiftedA_3__10_, 
        shiftedA_3__9_, shiftedA_3__8_, shiftedA_3__7_, shiftedA_3__6_, 
        shiftedA_3__5_, shiftedA_3__4_, shiftedA_3__3_, 1'b0, 1'b0, 1'b0}), 
        .b({n125, n125, n125, n125, n125, n125, n125, n125, n125, n125, n125, 
        n125, n125, n125, n125, n125, n125, n125, n125, n125, n125, n125, n125, 
        n125, n125, n125, n125, n125, n125, shiftedA_4__34_, shiftedA_4__33_, 
        shiftedA_4__32_, shiftedA_4__31_, shiftedA_4__30_, shiftedA_4__29_, 
        shiftedA_4__28_, shiftedA_4__27_, shiftedA_4__26_, shiftedA_4__25_, 
        shiftedA_4__24_, shiftedA_4__23_, shiftedA_4__22_, shiftedA_4__21_, 
        shiftedA_4__20_, shiftedA_4__19_, shiftedA_4__18_, shiftedA_4__17_, 
        shiftedA_4__16_, shiftedA_4__15_, shiftedA_4__14_, shiftedA_4__13_, 
        shiftedA_4__12_, shiftedA_4__11_, shiftedA_4__10_, shiftedA_4__9_, 
        shiftedA_4__8_, shiftedA_4__7_, shiftedA_4__6_, shiftedA_4__5_, 
        shiftedA_4__4_, 1'b0, 1'b0, 1'b0, 1'b0}), .c({n124, n124, n124, n124, 
        n124, n124, n124, n124, n124, n124, n124, n124, n124, n124, n124, n124, 
        n124, n124, n124, n124, n124, n124, n124, n124, n124, n124, n124, n124, 
        shiftedA_5__35_, shiftedA_5__34_, shiftedA_5__33_, shiftedA_5__32_, 
        shiftedA_5__31_, shiftedA_5__30_, shiftedA_5__29_, shiftedA_5__28_, 
        shiftedA_5__27_, shiftedA_5__26_, shiftedA_5__25_, shiftedA_5__24_, 
        shiftedA_5__23_, shiftedA_5__22_, shiftedA_5__21_, shiftedA_5__20_, 
        shiftedA_5__19_, shiftedA_5__18_, shiftedA_5__17_, shiftedA_5__16_, 
        shiftedA_5__15_, shiftedA_5__14_, shiftedA_5__13_, shiftedA_5__12_, 
        shiftedA_5__11_, shiftedA_5__10_, shiftedA_5__9_, shiftedA_5__8_, 
        shiftedA_5__7_, shiftedA_5__6_, shiftedA_5__5_, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .result(adderResult_level1[127:64]), .carry(
        carry_level1[127:64]) );
  BWAdder_60 level1_2__adder ( .a({n122, n122, n122, n122, n122, n122, n122, 
        n122, n122, n122, n122, n122, n122, n122, n122, n122, n122, n122, n122, 
        n122, n122, n122, n122, n122, n122, n122, n122, shiftedA_6__36_, 
        shiftedA_6__35_, shiftedA_6__34_, shiftedA_6__33_, shiftedA_6__32_, 
        shiftedA_6__31_, shiftedA_6__30_, shiftedA_6__29_, shiftedA_6__28_, 
        shiftedA_6__27_, shiftedA_6__26_, shiftedA_6__25_, shiftedA_6__24_, 
        shiftedA_6__23_, shiftedA_6__22_, shiftedA_6__21_, shiftedA_6__20_, 
        shiftedA_6__19_, shiftedA_6__18_, shiftedA_6__17_, shiftedA_6__16_, 
        shiftedA_6__15_, shiftedA_6__14_, shiftedA_6__13_, shiftedA_6__12_, 
        shiftedA_6__11_, shiftedA_6__10_, shiftedA_6__9_, shiftedA_6__8_, 
        shiftedA_6__7_, shiftedA_6__6_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .b({n119, n119, n119, n119, n119, n119, n119, n119, n119, n119, n119, 
        n119, n119, n119, n119, n119, n119, n119, n119, n119, n119, n119, n119, 
        n119, n119, n119, shiftedA_7__37_, shiftedA_7__36_, shiftedA_7__35_, 
        shiftedA_7__34_, shiftedA_7__33_, shiftedA_7__32_, shiftedA_7__31_, 
        shiftedA_7__30_, shiftedA_7__29_, shiftedA_7__28_, shiftedA_7__27_, 
        shiftedA_7__26_, shiftedA_7__25_, shiftedA_7__24_, shiftedA_7__23_, 
        shiftedA_7__22_, shiftedA_7__21_, shiftedA_7__20_, shiftedA_7__19_, 
        shiftedA_7__18_, shiftedA_7__17_, shiftedA_7__16_, shiftedA_7__15_, 
        shiftedA_7__14_, shiftedA_7__13_, shiftedA_7__12_, shiftedA_7__11_, 
        shiftedA_7__10_, shiftedA_7__9_, shiftedA_7__8_, shiftedA_7__7_, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({n118, n118, n118, n118, n118, 
        n118, n118, n118, n118, n118, n118, n118, n118, n118, n118, n118, n118, 
        n118, n118, n118, n118, n118, n118, n118, n118, shiftedA_8__38_, 
        shiftedA_8__37_, shiftedA_8__36_, shiftedA_8__35_, shiftedA_8__34_, 
        shiftedA_8__33_, shiftedA_8__32_, shiftedA_8__31_, shiftedA_8__30_, 
        shiftedA_8__29_, shiftedA_8__28_, shiftedA_8__27_, shiftedA_8__26_, 
        shiftedA_8__25_, shiftedA_8__24_, shiftedA_8__23_, shiftedA_8__22_, 
        shiftedA_8__21_, shiftedA_8__20_, shiftedA_8__19_, shiftedA_8__18_, 
        shiftedA_8__17_, shiftedA_8__16_, shiftedA_8__15_, shiftedA_8__14_, 
        shiftedA_8__13_, shiftedA_8__12_, shiftedA_8__11_, shiftedA_8__10_, 
        shiftedA_8__9_, shiftedA_8__8_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .result(adderResult_level1[191:128]), .carry(
        carry_level1[191:128]) );
  BWAdder_59 level1_3__adder ( .a({n116, n116, n116, n116, n116, n116, n116, 
        n116, n116, n116, n116, n116, n116, n116, n116, n116, n116, n116, n116, 
        n116, n116, n116, n116, n116, shiftedA_9__39_, shiftedA_9__38_, 
        shiftedA_9__37_, shiftedA_9__36_, shiftedA_9__35_, shiftedA_9__34_, 
        shiftedA_9__33_, shiftedA_9__32_, shiftedA_9__31_, shiftedA_9__30_, 
        shiftedA_9__29_, shiftedA_9__28_, shiftedA_9__27_, shiftedA_9__26_, 
        shiftedA_9__25_, shiftedA_9__24_, shiftedA_9__23_, shiftedA_9__22_, 
        shiftedA_9__21_, shiftedA_9__20_, shiftedA_9__19_, shiftedA_9__18_, 
        shiftedA_9__17_, shiftedA_9__16_, shiftedA_9__15_, shiftedA_9__14_, 
        shiftedA_9__13_, shiftedA_9__12_, shiftedA_9__11_, shiftedA_9__10_, 
        shiftedA_9__9_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .b({n113, n113, n113, n113, n113, n113, n113, n113, n113, n113, n113, 
        n113, n113, n113, n113, n113, n113, n113, n113, n113, n113, n113, n113, 
        shiftedA_10__40_, shiftedA_10__39_, shiftedA_10__38_, shiftedA_10__37_, 
        shiftedA_10__36_, shiftedA_10__35_, shiftedA_10__34_, shiftedA_10__33_, 
        shiftedA_10__32_, shiftedA_10__31_, shiftedA_10__30_, shiftedA_10__29_, 
        shiftedA_10__28_, shiftedA_10__27_, shiftedA_10__26_, shiftedA_10__25_, 
        shiftedA_10__24_, shiftedA_10__23_, shiftedA_10__22_, shiftedA_10__21_, 
        shiftedA_10__20_, shiftedA_10__19_, shiftedA_10__18_, shiftedA_10__17_, 
        shiftedA_10__16_, shiftedA_10__15_, shiftedA_10__14_, shiftedA_10__13_, 
        shiftedA_10__12_, shiftedA_10__11_, shiftedA_10__10_, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({n112, n112, n112, n112, 
        n112, n112, n112, n112, n112, n112, n112, n112, n112, n112, n112, n112, 
        n112, n112, n112, n112, n112, n112, shiftedA_11__41_, shiftedA_11__40_, 
        shiftedA_11__39_, shiftedA_11__38_, shiftedA_11__37_, shiftedA_11__36_, 
        shiftedA_11__35_, shiftedA_11__34_, shiftedA_11__33_, shiftedA_11__32_, 
        shiftedA_11__31_, shiftedA_11__30_, shiftedA_11__29_, shiftedA_11__28_, 
        shiftedA_11__27_, shiftedA_11__26_, shiftedA_11__25_, shiftedA_11__24_, 
        shiftedA_11__23_, shiftedA_11__22_, shiftedA_11__21_, shiftedA_11__20_, 
        shiftedA_11__19_, shiftedA_11__18_, shiftedA_11__17_, shiftedA_11__16_, 
        shiftedA_11__15_, shiftedA_11__14_, shiftedA_11__13_, shiftedA_11__12_, 
        shiftedA_11__11_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .result(adderResult_level1[255:192]), .carry(
        carry_level1[255:192]) );
  BWAdder_58 level1_4__adder ( .a({n109, n109, n109, n109, n109, n109, n109, 
        n109, n109, n109, n109, n109, n109, n109, n109, n109, n109, n109, n109, 
        n109, n109, shiftedA_12__42_, shiftedA_12__41_, shiftedA_12__40_, 
        shiftedA_12__39_, shiftedA_12__38_, shiftedA_12__37_, shiftedA_12__36_, 
        shiftedA_12__35_, shiftedA_12__34_, shiftedA_12__33_, shiftedA_12__32_, 
        shiftedA_12__31_, shiftedA_12__30_, shiftedA_12__29_, shiftedA_12__28_, 
        shiftedA_12__27_, shiftedA_12__26_, shiftedA_12__25_, shiftedA_12__24_, 
        shiftedA_12__23_, shiftedA_12__22_, shiftedA_12__21_, shiftedA_12__20_, 
        shiftedA_12__19_, shiftedA_12__18_, shiftedA_12__17_, shiftedA_12__16_, 
        shiftedA_12__15_, shiftedA_12__14_, shiftedA_12__13_, shiftedA_12__12_, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n108, n108, n108, n108, n108, n108, n108, n108, n108, n108, n108, n108, 
        n108, n108, n108, n108, n108, n108, n108, n108, shiftedA_13__43_, 
        shiftedA_13__42_, shiftedA_13__41_, shiftedA_13__40_, shiftedA_13__39_, 
        shiftedA_13__38_, shiftedA_13__37_, shiftedA_13__36_, shiftedA_13__35_, 
        shiftedA_13__34_, shiftedA_13__33_, shiftedA_13__32_, shiftedA_13__31_, 
        shiftedA_13__30_, shiftedA_13__29_, shiftedA_13__28_, shiftedA_13__27_, 
        shiftedA_13__26_, shiftedA_13__25_, shiftedA_13__24_, shiftedA_13__23_, 
        shiftedA_13__22_, shiftedA_13__21_, shiftedA_13__20_, shiftedA_13__19_, 
        shiftedA_13__18_, shiftedA_13__17_, shiftedA_13__16_, shiftedA_13__15_, 
        shiftedA_13__14_, shiftedA_13__13_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({n105, n105, n105, n105, 
        n105, n105, n105, n105, n105, n105, n105, n105, n105, n105, n105, n105, 
        n105, n105, n105, shiftedA_14__44_, shiftedA_14__43_, shiftedA_14__42_, 
        shiftedA_14__41_, shiftedA_14__40_, shiftedA_14__39_, shiftedA_14__38_, 
        shiftedA_14__37_, shiftedA_14__36_, shiftedA_14__35_, shiftedA_14__34_, 
        shiftedA_14__33_, shiftedA_14__32_, shiftedA_14__31_, shiftedA_14__30_, 
        shiftedA_14__29_, shiftedA_14__28_, shiftedA_14__27_, shiftedA_14__26_, 
        shiftedA_14__25_, shiftedA_14__24_, shiftedA_14__23_, shiftedA_14__22_, 
        shiftedA_14__21_, shiftedA_14__20_, shiftedA_14__19_, shiftedA_14__18_, 
        shiftedA_14__17_, shiftedA_14__16_, shiftedA_14__15_, shiftedA_14__14_, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .result(adderResult_level1[319:256]), .carry(
        carry_level1[319:256]) );
  BWAdder_57 level1_5__adder ( .a({n103, n103, n103, n103, n103, n103, n103, 
        n103, n103, n103, n103, n103, n103, n103, n103, n103, n103, n103, 
        shiftedA_15__45_, shiftedA_15__44_, shiftedA_15__43_, shiftedA_15__42_, 
        shiftedA_15__41_, shiftedA_15__40_, shiftedA_15__39_, shiftedA_15__38_, 
        shiftedA_15__37_, shiftedA_15__36_, shiftedA_15__35_, shiftedA_15__34_, 
        shiftedA_15__33_, shiftedA_15__32_, shiftedA_15__31_, shiftedA_15__30_, 
        shiftedA_15__29_, shiftedA_15__28_, shiftedA_15__27_, shiftedA_15__26_, 
        shiftedA_15__25_, shiftedA_15__24_, shiftedA_15__23_, shiftedA_15__22_, 
        shiftedA_15__21_, shiftedA_15__20_, shiftedA_15__19_, shiftedA_15__18_, 
        shiftedA_15__17_, shiftedA_15__16_, shiftedA_15__15_, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n102, n102, n102, n102, n102, n102, n102, n102, n102, n102, n102, n102, 
        n102, n102, n102, n102, n102, shiftedA_16__46_, shiftedA_16__45_, 
        shiftedA_16__44_, shiftedA_16__43_, shiftedA_16__42_, shiftedA_16__41_, 
        shiftedA_16__40_, shiftedA_16__39_, shiftedA_16__38_, shiftedA_16__37_, 
        shiftedA_16__36_, shiftedA_16__35_, shiftedA_16__34_, shiftedA_16__33_, 
        shiftedA_16__32_, shiftedA_16__31_, shiftedA_16__30_, shiftedA_16__29_, 
        shiftedA_16__28_, shiftedA_16__27_, shiftedA_16__26_, shiftedA_16__25_, 
        shiftedA_16__24_, shiftedA_16__23_, shiftedA_16__22_, shiftedA_16__21_, 
        shiftedA_16__20_, shiftedA_16__19_, shiftedA_16__18_, shiftedA_16__17_, 
        shiftedA_16__16_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({n99, n99, n99, n99, 
        n99, n99, n99, n99, n99, n99, n99, n99, n99, n99, n99, n99, 
        shiftedA_17__47_, shiftedA_17__46_, shiftedA_17__45_, shiftedA_17__44_, 
        shiftedA_17__43_, shiftedA_17__42_, shiftedA_17__41_, shiftedA_17__40_, 
        shiftedA_17__39_, shiftedA_17__38_, shiftedA_17__37_, shiftedA_17__36_, 
        shiftedA_17__35_, shiftedA_17__34_, shiftedA_17__33_, shiftedA_17__32_, 
        shiftedA_17__31_, shiftedA_17__30_, shiftedA_17__29_, shiftedA_17__28_, 
        shiftedA_17__27_, shiftedA_17__26_, shiftedA_17__25_, shiftedA_17__24_, 
        shiftedA_17__23_, shiftedA_17__22_, shiftedA_17__21_, shiftedA_17__20_, 
        shiftedA_17__19_, shiftedA_17__18_, shiftedA_17__17_, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .result(adderResult_level1[383:320]), .carry(
        carry_level1[383:320]) );
  BWAdder_56 level1_6__adder ( .a({shiftedA_18__63_, shiftedA_18__63_, 
        shiftedA_18__63_, shiftedA_18__63_, shiftedA_18__63_, shiftedA_18__63_, 
        shiftedA_18__63_, shiftedA_18__63_, shiftedA_18__63_, shiftedA_18__63_, 
        shiftedA_18__63_, shiftedA_18__63_, shiftedA_18__63_, shiftedA_18__63_, 
        shiftedA_18__63_, shiftedA_18__48_, shiftedA_18__47_, shiftedA_18__46_, 
        shiftedA_18__45_, shiftedA_18__44_, shiftedA_18__43_, shiftedA_18__42_, 
        shiftedA_18__41_, shiftedA_18__40_, shiftedA_18__39_, shiftedA_18__38_, 
        shiftedA_18__37_, shiftedA_18__36_, shiftedA_18__35_, shiftedA_18__34_, 
        shiftedA_18__33_, shiftedA_18__32_, shiftedA_18__31_, shiftedA_18__30_, 
        shiftedA_18__29_, shiftedA_18__28_, shiftedA_18__27_, shiftedA_18__26_, 
        shiftedA_18__25_, shiftedA_18__24_, shiftedA_18__23_, shiftedA_18__22_, 
        shiftedA_18__21_, shiftedA_18__20_, shiftedA_18__19_, shiftedA_18__18_, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_19__63_, 
        shiftedA_19__63_, shiftedA_19__63_, shiftedA_19__63_, shiftedA_19__63_, 
        shiftedA_19__63_, shiftedA_19__63_, shiftedA_19__63_, shiftedA_19__63_, 
        shiftedA_19__63_, shiftedA_19__63_, shiftedA_19__63_, shiftedA_19__63_, 
        shiftedA_19__63_, shiftedA_19__49_, shiftedA_19__48_, shiftedA_19__47_, 
        shiftedA_19__46_, shiftedA_19__45_, shiftedA_19__44_, shiftedA_19__43_, 
        shiftedA_19__42_, shiftedA_19__41_, shiftedA_19__40_, shiftedA_19__39_, 
        shiftedA_19__38_, shiftedA_19__37_, shiftedA_19__36_, shiftedA_19__35_, 
        shiftedA_19__34_, shiftedA_19__33_, shiftedA_19__32_, shiftedA_19__31_, 
        shiftedA_19__30_, shiftedA_19__29_, shiftedA_19__28_, shiftedA_19__27_, 
        shiftedA_19__26_, shiftedA_19__25_, shiftedA_19__24_, shiftedA_19__23_, 
        shiftedA_19__22_, shiftedA_19__21_, shiftedA_19__20_, shiftedA_19__19_, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_20__63_, 
        shiftedA_20__63_, shiftedA_20__63_, shiftedA_20__63_, shiftedA_20__63_, 
        shiftedA_20__63_, shiftedA_20__63_, shiftedA_20__63_, shiftedA_20__63_, 
        shiftedA_20__63_, shiftedA_20__63_, shiftedA_20__63_, shiftedA_20__63_, 
        shiftedA_20__50_, shiftedA_20__49_, shiftedA_20__48_, shiftedA_20__47_, 
        shiftedA_20__46_, shiftedA_20__45_, shiftedA_20__44_, shiftedA_20__43_, 
        shiftedA_20__42_, shiftedA_20__41_, shiftedA_20__40_, shiftedA_20__39_, 
        shiftedA_20__38_, shiftedA_20__37_, shiftedA_20__36_, shiftedA_20__35_, 
        shiftedA_20__34_, shiftedA_20__33_, shiftedA_20__32_, shiftedA_20__31_, 
        shiftedA_20__30_, shiftedA_20__29_, shiftedA_20__28_, shiftedA_20__27_, 
        shiftedA_20__26_, shiftedA_20__25_, shiftedA_20__24_, shiftedA_20__23_, 
        shiftedA_20__22_, shiftedA_20__21_, shiftedA_20__20_, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(adderResult_level1[447:384]), 
        .carry(carry_level1[447:384]) );
  BWAdder_55 level1_7__adder ( .a({shiftedA_21__63_, shiftedA_21__63_, 
        shiftedA_21__63_, shiftedA_21__63_, shiftedA_21__63_, shiftedA_21__63_, 
        shiftedA_21__63_, shiftedA_21__63_, shiftedA_21__63_, shiftedA_21__63_, 
        shiftedA_21__63_, shiftedA_21__63_, shiftedA_21__51_, shiftedA_21__50_, 
        shiftedA_21__49_, shiftedA_21__48_, shiftedA_21__47_, shiftedA_21__46_, 
        shiftedA_21__45_, shiftedA_21__44_, shiftedA_21__43_, shiftedA_21__42_, 
        shiftedA_21__41_, shiftedA_21__40_, shiftedA_21__39_, shiftedA_21__38_, 
        shiftedA_21__37_, shiftedA_21__36_, shiftedA_21__35_, shiftedA_21__34_, 
        shiftedA_21__33_, shiftedA_21__32_, shiftedA_21__31_, shiftedA_21__30_, 
        shiftedA_21__29_, shiftedA_21__28_, shiftedA_21__27_, shiftedA_21__26_, 
        shiftedA_21__25_, shiftedA_21__24_, shiftedA_21__23_, shiftedA_21__22_, 
        shiftedA_21__21_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_22__63_, shiftedA_22__63_, shiftedA_22__63_, shiftedA_22__63_, 
        shiftedA_22__63_, shiftedA_22__63_, shiftedA_22__63_, shiftedA_22__63_, 
        shiftedA_22__63_, shiftedA_22__63_, shiftedA_22__63_, shiftedA_22__52_, 
        shiftedA_22__51_, shiftedA_22__50_, shiftedA_22__49_, shiftedA_22__48_, 
        shiftedA_22__47_, shiftedA_22__46_, shiftedA_22__45_, shiftedA_22__44_, 
        shiftedA_22__43_, shiftedA_22__42_, shiftedA_22__41_, shiftedA_22__40_, 
        shiftedA_22__39_, shiftedA_22__38_, shiftedA_22__37_, shiftedA_22__36_, 
        shiftedA_22__35_, shiftedA_22__34_, shiftedA_22__33_, shiftedA_22__32_, 
        shiftedA_22__31_, shiftedA_22__30_, shiftedA_22__29_, shiftedA_22__28_, 
        shiftedA_22__27_, shiftedA_22__26_, shiftedA_22__25_, shiftedA_22__24_, 
        shiftedA_22__23_, shiftedA_22__22_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_23__63_, shiftedA_23__63_, 
        shiftedA_23__63_, shiftedA_23__63_, shiftedA_23__63_, shiftedA_23__63_, 
        shiftedA_23__63_, shiftedA_23__63_, shiftedA_23__63_, shiftedA_23__63_, 
        shiftedA_23__53_, shiftedA_23__52_, shiftedA_23__51_, shiftedA_23__50_, 
        shiftedA_23__49_, shiftedA_23__48_, shiftedA_23__47_, shiftedA_23__46_, 
        shiftedA_23__45_, shiftedA_23__44_, shiftedA_23__43_, shiftedA_23__42_, 
        shiftedA_23__41_, shiftedA_23__40_, shiftedA_23__39_, shiftedA_23__38_, 
        shiftedA_23__37_, shiftedA_23__36_, shiftedA_23__35_, shiftedA_23__34_, 
        shiftedA_23__33_, shiftedA_23__32_, shiftedA_23__31_, shiftedA_23__30_, 
        shiftedA_23__29_, shiftedA_23__28_, shiftedA_23__27_, shiftedA_23__26_, 
        shiftedA_23__25_, shiftedA_23__24_, shiftedA_23__23_, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[511:448]), .carry(carry_level1[511:448]) );
  BWAdder_54 level1_8__adder ( .a({shiftedA_24__63_, shiftedA_24__63_, 
        shiftedA_24__63_, shiftedA_24__63_, shiftedA_24__63_, shiftedA_24__63_, 
        shiftedA_24__63_, shiftedA_24__63_, shiftedA_24__63_, shiftedA_24__54_, 
        shiftedA_24__53_, shiftedA_24__52_, shiftedA_24__51_, shiftedA_24__50_, 
        shiftedA_24__49_, shiftedA_24__48_, shiftedA_24__47_, shiftedA_24__46_, 
        shiftedA_24__45_, shiftedA_24__44_, shiftedA_24__43_, shiftedA_24__42_, 
        shiftedA_24__41_, shiftedA_24__40_, shiftedA_24__39_, shiftedA_24__38_, 
        shiftedA_24__37_, shiftedA_24__36_, shiftedA_24__35_, shiftedA_24__34_, 
        shiftedA_24__33_, shiftedA_24__32_, shiftedA_24__31_, shiftedA_24__30_, 
        shiftedA_24__29_, shiftedA_24__28_, shiftedA_24__27_, shiftedA_24__26_, 
        shiftedA_24__25_, shiftedA_24__24_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_25__63_, 
        shiftedA_25__63_, shiftedA_25__63_, shiftedA_25__63_, shiftedA_25__63_, 
        shiftedA_25__63_, shiftedA_25__63_, shiftedA_25__63_, shiftedA_25__55_, 
        shiftedA_25__54_, shiftedA_25__53_, shiftedA_25__52_, shiftedA_25__51_, 
        shiftedA_25__50_, shiftedA_25__49_, shiftedA_25__48_, shiftedA_25__47_, 
        shiftedA_25__46_, shiftedA_25__45_, shiftedA_25__44_, shiftedA_25__43_, 
        shiftedA_25__42_, shiftedA_25__41_, shiftedA_25__40_, shiftedA_25__39_, 
        shiftedA_25__38_, shiftedA_25__37_, shiftedA_25__36_, shiftedA_25__35_, 
        shiftedA_25__34_, shiftedA_25__33_, shiftedA_25__32_, shiftedA_25__31_, 
        shiftedA_25__30_, shiftedA_25__29_, shiftedA_25__28_, shiftedA_25__27_, 
        shiftedA_25__26_, shiftedA_25__25_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_26__63_, 
        shiftedA_26__63_, shiftedA_26__63_, shiftedA_26__63_, shiftedA_26__63_, 
        shiftedA_26__63_, shiftedA_26__63_, shiftedA_26__56_, shiftedA_26__55_, 
        shiftedA_26__54_, shiftedA_26__53_, shiftedA_26__52_, shiftedA_26__51_, 
        shiftedA_26__50_, shiftedA_26__49_, shiftedA_26__48_, shiftedA_26__47_, 
        shiftedA_26__46_, shiftedA_26__45_, shiftedA_26__44_, shiftedA_26__43_, 
        shiftedA_26__42_, shiftedA_26__41_, shiftedA_26__40_, shiftedA_26__39_, 
        shiftedA_26__38_, shiftedA_26__37_, shiftedA_26__36_, shiftedA_26__35_, 
        shiftedA_26__34_, shiftedA_26__33_, shiftedA_26__32_, shiftedA_26__31_, 
        shiftedA_26__30_, shiftedA_26__29_, shiftedA_26__28_, shiftedA_26__27_, 
        shiftedA_26__26_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(adderResult_level1[575:512]), 
        .carry(carry_level1[575:512]) );
  BWAdder_53 level1_9__adder ( .a({shiftedA_27__63_, shiftedA_27__63_, 
        shiftedA_27__63_, shiftedA_27__63_, shiftedA_27__63_, shiftedA_27__63_, 
        shiftedA_27__57_, shiftedA_27__56_, shiftedA_27__55_, shiftedA_27__54_, 
        shiftedA_27__53_, shiftedA_27__52_, shiftedA_27__51_, shiftedA_27__50_, 
        shiftedA_27__49_, shiftedA_27__48_, shiftedA_27__47_, shiftedA_27__46_, 
        shiftedA_27__45_, shiftedA_27__44_, shiftedA_27__43_, shiftedA_27__42_, 
        shiftedA_27__41_, shiftedA_27__40_, shiftedA_27__39_, shiftedA_27__38_, 
        shiftedA_27__37_, shiftedA_27__36_, shiftedA_27__35_, shiftedA_27__34_, 
        shiftedA_27__33_, shiftedA_27__32_, shiftedA_27__31_, shiftedA_27__30_, 
        shiftedA_27__29_, shiftedA_27__28_, shiftedA_27__27_, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_28__63_, shiftedA_28__63_, shiftedA_28__63_, shiftedA_28__63_, 
        shiftedA_28__63_, shiftedA_28__58_, shiftedA_28__57_, shiftedA_28__56_, 
        shiftedA_28__55_, shiftedA_28__54_, shiftedA_28__53_, shiftedA_28__52_, 
        shiftedA_28__51_, shiftedA_28__50_, shiftedA_28__49_, shiftedA_28__48_, 
        shiftedA_28__47_, shiftedA_28__46_, shiftedA_28__45_, shiftedA_28__44_, 
        shiftedA_28__43_, shiftedA_28__42_, shiftedA_28__41_, shiftedA_28__40_, 
        shiftedA_28__39_, shiftedA_28__38_, shiftedA_28__37_, shiftedA_28__36_, 
        shiftedA_28__35_, shiftedA_28__34_, shiftedA_28__33_, shiftedA_28__32_, 
        shiftedA_28__31_, shiftedA_28__30_, shiftedA_28__29_, shiftedA_28__28_, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_29__63_, shiftedA_29__63_, 
        shiftedA_29__63_, shiftedA_29__63_, shiftedA_29__59_, shiftedA_29__58_, 
        shiftedA_29__57_, shiftedA_29__56_, shiftedA_29__55_, shiftedA_29__54_, 
        shiftedA_29__53_, shiftedA_29__52_, shiftedA_29__51_, shiftedA_29__50_, 
        shiftedA_29__49_, shiftedA_29__48_, shiftedA_29__47_, shiftedA_29__46_, 
        shiftedA_29__45_, shiftedA_29__44_, shiftedA_29__43_, shiftedA_29__42_, 
        shiftedA_29__41_, shiftedA_29__40_, shiftedA_29__39_, shiftedA_29__38_, 
        shiftedA_29__37_, shiftedA_29__36_, shiftedA_29__35_, shiftedA_29__34_, 
        shiftedA_29__33_, shiftedA_29__32_, shiftedA_29__31_, shiftedA_29__30_, 
        shiftedA_29__29_, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[639:576]), .carry(carry_level1[639:576]) );
  BWAdder_52 level1_10__adder ( .a({shiftedA_30__63_, shiftedA_30__63_, 
        shiftedA_30__63_, shiftedA_30__60_, shiftedA_30__59_, shiftedA_30__58_, 
        shiftedA_30__57_, shiftedA_30__56_, shiftedA_30__55_, shiftedA_30__54_, 
        shiftedA_30__53_, shiftedA_30__52_, shiftedA_30__51_, shiftedA_30__50_, 
        shiftedA_30__49_, shiftedA_30__48_, shiftedA_30__47_, shiftedA_30__46_, 
        shiftedA_30__45_, shiftedA_30__44_, shiftedA_30__43_, shiftedA_30__42_, 
        shiftedA_30__41_, shiftedA_30__40_, shiftedA_30__39_, shiftedA_30__38_, 
        shiftedA_30__37_, shiftedA_30__36_, shiftedA_30__35_, shiftedA_30__34_, 
        shiftedA_30__33_, shiftedA_30__32_, shiftedA_30__31_, shiftedA_30__30_, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_32__63_, 
        shiftedA_32__63_, shiftedA_33__63_, shiftedA_34__63_, shiftedA_35__63_, 
        shiftedA_36__63_, shiftedA_37__63_, shiftedA_38__63_, shiftedA_39__63_, 
        shiftedA_40__63_, shiftedA_41__63_, shiftedA_42__63_, shiftedA_43__63_, 
        shiftedA_44__63_, shiftedA_45__63_, n100, n101, n104, n106, n107, n110, 
        n111, n114, n115, n117, n120, n121, n123, n126, n127, n129, n132, n133, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_32__63_, 
        shiftedA_33__63_, shiftedA_34__63_, shiftedA_35__63_, shiftedA_36__63_, 
        shiftedA_37__63_, shiftedA_38__63_, shiftedA_39__63_, shiftedA_40__63_, 
        shiftedA_41__63_, shiftedA_42__63_, shiftedA_43__63_, shiftedA_44__63_, 
        shiftedA_45__63_, n100, n101, n104, n106, n107, n110, n111, n114, n115, 
        n117, n120, n121, n123, n126, n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(adderResult_level1[703:640]), 
        .carry(carry_level1[703:640]) );
  BWAdder_51 level1_11__adder ( .a({shiftedA_33__63_, shiftedA_34__63_, 
        shiftedA_35__63_, shiftedA_36__63_, shiftedA_37__63_, shiftedA_38__63_, 
        shiftedA_39__63_, shiftedA_40__63_, shiftedA_41__63_, shiftedA_42__63_, 
        shiftedA_43__63_, shiftedA_44__63_, shiftedA_45__63_, n100, n101, n104, 
        n106, n107, n110, n111, n114, n115, n117, n120, n121, n123, n126, n127, 
        n129, n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_34__63_, shiftedA_35__63_, shiftedA_36__63_, shiftedA_37__63_, 
        shiftedA_38__63_, shiftedA_39__63_, shiftedA_40__63_, shiftedA_41__63_, 
        shiftedA_42__63_, shiftedA_43__63_, shiftedA_44__63_, shiftedA_45__63_, 
        n100, n101, n104, n106, n107, n110, n111, n114, n115, n117, n120, n121, 
        n123, n126, n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_35__63_, shiftedA_36__63_, 
        shiftedA_37__63_, shiftedA_38__63_, shiftedA_39__63_, shiftedA_40__63_, 
        shiftedA_41__63_, shiftedA_42__63_, shiftedA_43__63_, shiftedA_44__63_, 
        shiftedA_45__63_, n100, n101, n104, n106, n107, n110, n111, n114, n115, 
        n117, n120, n121, n123, n126, n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[767:704]), .carry(carry_level1[767:704]) );
  BWAdder_50 level1_12__adder ( .a({shiftedA_36__63_, shiftedA_37__63_, 
        shiftedA_38__63_, shiftedA_39__63_, shiftedA_40__63_, shiftedA_41__63_, 
        shiftedA_42__63_, shiftedA_43__63_, shiftedA_44__63_, shiftedA_45__63_, 
        n100, n101, n104, n106, n107, n110, n111, n114, n115, n117, n120, n121, 
        n123, n126, n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_37__63_, 
        shiftedA_38__63_, shiftedA_39__63_, shiftedA_40__63_, shiftedA_41__63_, 
        shiftedA_42__63_, shiftedA_43__63_, shiftedA_44__63_, shiftedA_45__63_, 
        n100, n101, n104, n106, n107, n110, n111, n114, n115, n117, n120, n121, 
        n123, n126, n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_38__63_, 
        shiftedA_39__63_, shiftedA_40__63_, shiftedA_41__63_, shiftedA_42__63_, 
        shiftedA_43__63_, shiftedA_44__63_, shiftedA_45__63_, n100, n101, n104, 
        n106, n107, n110, n111, n114, n115, n117, n120, n121, n123, n126, n127, 
        n129, n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(adderResult_level1[831:768]), 
        .carry(carry_level1[831:768]) );
  BWAdder_49 level1_13__adder ( .a({shiftedA_39__63_, shiftedA_40__63_, 
        shiftedA_41__63_, shiftedA_42__63_, shiftedA_43__63_, shiftedA_44__63_, 
        shiftedA_45__63_, n100, n101, n104, n106, n107, n110, n111, n114, n115, 
        n117, n120, n121, n123, n126, n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_40__63_, shiftedA_41__63_, shiftedA_42__63_, shiftedA_43__63_, 
        shiftedA_44__63_, shiftedA_45__63_, n100, n101, n104, n106, n107, n110, 
        n111, n114, n115, n117, n120, n121, n123, n126, n127, n129, n132, n133, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_41__63_, shiftedA_42__63_, 
        shiftedA_43__63_, shiftedA_44__63_, shiftedA_45__63_, n100, n101, n104, 
        n106, n107, n110, n111, n114, n115, n117, n120, n121, n123, n126, n127, 
        n129, n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[895:832]), .carry(carry_level1[895:832]) );
  BWAdder_48 level1_14__adder ( .a({shiftedA_42__63_, shiftedA_43__63_, 
        shiftedA_44__63_, shiftedA_45__63_, n100, n101, n104, n106, n107, n110, 
        n111, n114, n115, n117, n120, n121, n123, n126, n127, n129, n132, n133, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({shiftedA_43__63_, 
        shiftedA_44__63_, shiftedA_45__63_, n100, n101, n104, n106, n107, n110, 
        n111, n114, n115, n117, n120, n121, n123, n126, n127, n129, n132, n133, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({shiftedA_44__63_, 
        shiftedA_45__63_, n100, n101, n104, n106, n107, n110, n111, n114, n115, 
        n117, n120, n121, n123, n126, n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(adderResult_level1[959:896]), 
        .carry(carry_level1[959:896]) );
  BWAdder_47 level1_15__adder ( .a({shiftedA_45__63_, n100, n101, n104, n106, 
        n107, n110, n111, n114, n115, n117, n120, n121, n123, n126, n127, n129, 
        n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .b({n100, n101, n104, n106, n107, n110, n111, n114, n115, n117, n120, 
        n121, n123, n126, n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .c({n101, n104, n106, n107, n110, n111, 
        n114, n115, n117, n120, n121, n123, n126, n127, n129, n132, n133, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[1023:960]), .carry(carry_level1[1023:960]) );
  BWAdder_46 level1_16__adder ( .a({n104, n106, n107, n110, n111, n114, n115, 
        n117, n120, n121, n123, n126, n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n106, n107, 
        n110, n111, n114, n115, n117, n120, n121, n123, n126, n127, n129, n132, 
        n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .c({n107, n110, n111, n114, n115, n117, n120, n121, n123, 
        n126, n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[1087:1024]), .carry(carry_level1[1087:1024]) );
  BWAdder_45 level1_17__adder ( .a({n110, n111, n114, n115, n117, n120, n121, 
        n123, n126, n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n111, n114, 
        n115, n117, n120, n121, n123, n126, n127, n129, n132, n133, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .c({n114, n115, n117, n120, n121, n123, n126, n127, n129, 
        n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[1151:1088]), .carry(carry_level1[1151:1088]) );
  BWAdder_44 level1_18__adder ( .a({n115, n117, n120, n121, n123, n126, n127, 
        n129, n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n117, n120, 
        n121, n123, n126, n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .c({n120, n121, n123, n126, n127, n129, n132, n133, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[1215:1152]), .carry(carry_level1[1215:1152]) );
  BWAdder_43 level1_19__adder ( .a({n121, n123, n126, n127, n129, n132, n133, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n123, n126, 
        n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .c({n126, n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[1279:1216]), .carry(carry_level1[1279:1216]) );
  BWAdder_42 level1_20__adder ( .a({n127, n129, n132, n133, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({n129, n132, 
        n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .c({n132, n133, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .result(
        adderResult_level1[1343:1280]), .carry(carry_level1[1343:1280]) );
  BWAdder_41 level2_a_0__adder ( .a(adderResult_level1[63:0]), .b(
        adderResult_level1[127:64]), .c(adderResult_level1[191:128]), .result(
        adderResult_level2[63:0]), .carry(carry_level2[63:0]) );
  BWAdder_40 level2_a_1__adder ( .a(adderResult_level1[255:192]), .b(
        adderResult_level1[319:256]), .c(adderResult_level1[383:320]), 
        .result(adderResult_level2[127:64]), .carry(carry_level2[127:64]) );
  BWAdder_39 level2_a_2__adder ( .a(adderResult_level1[447:384]), .b(
        adderResult_level1[511:448]), .c(adderResult_level1[575:512]), 
        .result(adderResult_level2[191:128]), .carry(carry_level2[191:128]) );
  BWAdder_38 level2_a_3__adder ( .a(adderResult_level1[639:576]), .b(
        adderResult_level1[703:640]), .c(adderResult_level1[767:704]), 
        .result(adderResult_level2[255:192]), .carry(carry_level2[255:192]) );
  BWAdder_37 level2_a_4__adder ( .a(adderResult_level1[831:768]), .b(
        adderResult_level1[895:832]), .c(adderResult_level1[959:896]), 
        .result(adderResult_level2[319:256]), .carry(carry_level2[319:256]) );
  BWAdder_36 level2_a_5__adder ( .a(adderResult_level1[1023:960]), .b(
        adderResult_level1[1087:1024]), .c(adderResult_level1[1151:1088]), 
        .result(adderResult_level2[383:320]), .carry(carry_level2[383:320]) );
  BWAdder_35 level2_a_6__adder ( .a(adderResult_level1[1215:1152]), .b(
        adderResult_level1[1279:1216]), .c(adderResult_level1[1343:1280]), 
        .result(adderResult_level2[447:384]), .carry(carry_level2[447:384]) );
  BWAdder_34 level2_b_0__adder ( .a({carry_level1[63:1], 1'b0}), .b({
        carry_level1[127:65], 1'b0}), .c({carry_level1[191:129], 1'b0}), 
        .result(adderResult_level2[511:448]), .carry(carry_level2[511:448]) );
  BWAdder_33 level2_b_1__adder ( .a({carry_level1[255:193], 1'b0}), .b({
        carry_level1[319:257], 1'b0}), .c({carry_level1[383:321], 1'b0}), 
        .result(adderResult_level2[575:512]), .carry(carry_level2[575:512]) );
  BWAdder_32 level2_b_2__adder ( .a({carry_level1[447:385], 1'b0}), .b({
        carry_level1[511:449], 1'b0}), .c({carry_level1[575:513], 1'b0}), 
        .result(adderResult_level2[639:576]), .carry(carry_level2[639:576]) );
  BWAdder_31 level2_b_3__adder ( .a({carry_level1[639:577], 1'b0}), .b({
        carry_level1[703:641], 1'b0}), .c({carry_level1[767:705], 1'b0}), 
        .result(adderResult_level2[703:640]), .carry(carry_level2[703:640]) );
  BWAdder_30 level2_b_4__adder ( .a({carry_level1[831:769], 1'b0}), .b({
        carry_level1[895:833], 1'b0}), .c({carry_level1[959:897], 1'b0}), 
        .result(adderResult_level2[767:704]), .carry(carry_level2[767:704]) );
  BWAdder_29 level2_b_5__adder ( .a({carry_level1[1023:961], 1'b0}), .b({
        carry_level1[1087:1025], 1'b0}), .c({carry_level1[1151:1089], 1'b0}), 
        .result(adderResult_level2[831:768]), .carry(carry_level2[831:768]) );
  BWAdder_28 level2_b_6__adder ( .a({carry_level1[1215:1153], 1'b0}), .b({
        carry_level1[1279:1217], 1'b0}), .c({carry_level1[1343:1281], 1'b0}), 
        .result(adderResult_level2[895:832]), .carry(carry_level2[895:832]) );
  BWAdder_27 level3_a_0__adder ( .a(adderResult_level2[63:0]), .b(
        adderResult_level2[127:64]), .c(adderResult_level2[191:128]), .result(
        adderResult_level3[63:0]), .carry(carry_level3[63:0]) );
  BWAdder_26 level3_a_1__adder ( .a(adderResult_level2[255:192]), .b(
        adderResult_level2[319:256]), .c(adderResult_level2[383:320]), 
        .result(adderResult_level3[127:64]), .carry(carry_level3[127:64]) );
  BWAdder_25 level3_a_2__adder ( .a(adderResult_level2[447:384]), .b(
        adderResult_level2[511:448]), .c(adderResult_level2[575:512]), 
        .result(adderResult_level3[191:128]), .carry(carry_level3[191:128]) );
  BWAdder_24 level3_a_3__adder ( .a(adderResult_level2[639:576]), .b(
        adderResult_level2[703:640]), .c(adderResult_level2[767:704]), 
        .result(adderResult_level3[255:192]), .carry(carry_level3[255:192]) );
  BWAdder_23 level3_b_0__adder ( .a({carry_level2[63:1], 1'b0}), .b({
        carry_level2[127:65], 1'b0}), .c({carry_level2[191:129], 1'b0}), 
        .result(adderResult_level3[319:256]), .carry(carry_level3[319:256]) );
  BWAdder_22 level3_b_1__adder ( .a({carry_level2[255:193], 1'b0}), .b({
        carry_level2[319:257], 1'b0}), .c({carry_level2[383:321], 1'b0}), 
        .result(adderResult_level3[383:320]), .carry(carry_level3[383:320]) );
  BWAdder_21 level3_b_2__adder ( .a({carry_level2[447:385], 1'b0}), .b({
        carry_level2[511:449], 1'b0}), .c({carry_level2[575:513], 1'b0}), 
        .result(adderResult_level3[447:384]), .carry(carry_level3[447:384]) );
  BWAdder_20 level3_b_3__adder ( .a({carry_level2[639:577], 1'b0}), .b({
        carry_level2[703:641], 1'b0}), .c({carry_level2[767:705], 1'b0}), 
        .result(adderResult_level3[511:448]), .carry(carry_level3[511:448]) );
  BWAdder_19 adder ( .a(adderResult_level2[831:768]), .b(
        adderResult_level2[895:832]), .c({carry_level2[831:769], 1'b0}), 
        .result(adderResult_level3[575:512]), .carry(carry_level3[575:512]) );
  BWAdder_18 level4_a_0__adder ( .a(adderResult_level3[63:0]), .b(
        adderResult_level3[127:64]), .c(adderResult_level3[191:128]), .result(
        adderResult_level4[63:0]), .carry(carry_level4[63:0]) );
  BWAdder_17 level4_a_1__adder ( .a(adderResult_level3[255:192]), .b(
        adderResult_level3[319:256]), .c(adderResult_level3[383:320]), 
        .result(adderResult_level4[127:64]), .carry(carry_level4[127:64]) );
  BWAdder_16 level4_a_2__adder ( .a(adderResult_level3[447:384]), .b(
        adderResult_level3[511:448]), .c(adderResult_level3[575:512]), 
        .result(adderResult_level4[191:128]), .carry(carry_level4[191:128]) );
  BWAdder_15 level4_b_0__adder ( .a({carry_level3[63:1], 1'b0}), .b({
        carry_level3[127:65], 1'b0}), .c({carry_level3[191:129], 1'b0}), 
        .result(adderResult_level4[255:192]), .carry(carry_level4[255:192]) );
  BWAdder_14 level4_b_1__adder ( .a({carry_level3[255:193], 1'b0}), .b({
        carry_level3[319:257], 1'b0}), .c({carry_level3[383:321], 1'b0}), 
        .result(adderResult_level4[319:256]), .carry(carry_level4[319:256]) );
  BWAdder_13 level4_b_2__adder ( .a({carry_level3[447:385], 1'b0}), .b({
        carry_level3[511:449], 1'b0}), .c({carry_level3[575:513], 1'b0}), 
        .result(adderResult_level4[383:320]), .carry(carry_level4[383:320]) );
  BWAdder_12 level5_a_0__adder ( .a(adderResult_level4[63:0]), .b(
        adderResult_level4[127:64]), .c(adderResult_level4[191:128]), .result(
        adderResult_level5[63:0]), .carry(carry_level5[63:0]) );
  BWAdder_11 level5_a_1__adder ( .a(adderResult_level4[255:192]), .b(
        adderResult_level4[319:256]), .c(adderResult_level4[383:320]), 
        .result(adderResult_level5[127:64]), .carry(carry_level5[127:64]) );
  BWAdder_10 level5_b_0__adder ( .a({carry_level4[63:1], 1'b0}), .b({
        carry_level4[127:65], 1'b0}), .c({carry_level4[191:129], 1'b0}), 
        .result(adderResult_level5[191:128]), .carry(carry_level5[191:128]) );
  BWAdder_9 level5_b_1__adder ( .a({carry_level4[255:193], 1'b0}), .b({
        carry_level4[319:257], 1'b0}), .c({carry_level4[383:321], 1'b0}), 
        .result(adderResult_level5[255:192]), .carry(carry_level5[255:192]) );
  BWAdder_8 adder_0 ( .a(adderResult_level5[63:0]), .b(
        adderResult_level5[127:64]), .c(adderResult_level5[191:128]), .result(
        adderResult_level6[63:0]), .carry(carry_level6[63:0]) );
  BWAdder_7 adder_1 ( .a(adderResult_level5[255:192]), .b({carry_level5[63:1], 
        1'b0}), .c({carry_level5[127:65], 1'b0}), .result(
        adderResult_level6[127:64]), .carry(carry_level6[127:64]) );
  BWAdder_6 adder_2 ( .a({carry_level5[191:129], 1'b0}), .b({
        carry_level5[255:193], 1'b0}), .c({carry_level2[895:833], 1'b0}), 
        .result(adderResult_level6[191:128]), .carry(carry_level6[191:128]) );
  BWAdder_5 adder_3 ( .a(adderResult_level6[63:0]), .b(
        adderResult_level6[127:64]), .c(adderResult_level6[191:128]), .result(
        adderResult_level7[63:0]), .carry(carry_level7[63:0]) );
  BWAdder_4 adder_4 ( .a({carry_level6[63:1], 1'b0}), .b({carry_level6[127:65], 
        1'b0}), .c({carry_level6[191:129], 1'b0}), .result(
        adderResult_level7[127:64]), .carry(carry_level7[127:64]) );
  BWAdder_3 adder_5 ( .a(adderResult_level7[63:0]), .b(
        adderResult_level7[127:64]), .c({carry_level7[63:1], 1'b0}), .result(
        adderResult_level8), .carry(carry_level8) );
  BWAdder_2 adder_6 ( .a(adderResult_level8), .b({carry_level7[127:65], 1'b0}), 
        .c({carry_level8[63:1], 1'b0}), .result(adderResult_level9), .carry(
        carry_level9) );
  BWAdder_1 adder_7 ( .a(adderResult_level9), .b({n133, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .c({carry_level9[63:1], 1'b0}), .result(adderResult_level10), .carry(
        carry_level10) );
  CRAdder_64 CRAdd ( .a(adderResult_level10), .b({carry_level10[63:1], 1'b0}), 
        .cin(1'b0), .sum(result) );
  OR2_X1 U1089 ( .A1(n159), .A2(n172), .ZN(n63) );
  OR2_X1 U1090 ( .A1(n158), .A2(n172), .ZN(n64) );
  OR2_X1 U1091 ( .A1(n138), .A2(n197), .ZN(n65) );
  OR2_X1 U1092 ( .A1(n157), .A2(n172), .ZN(n66) );
  OR2_X1 U1093 ( .A1(n138), .A2(n196), .ZN(n67) );
  OR2_X1 U1094 ( .A1(n138), .A2(n195), .ZN(n68) );
  OR2_X1 U1095 ( .A1(n156), .A2(n172), .ZN(n69) );
  OR2_X1 U1096 ( .A1(n155), .A2(n172), .ZN(n70) );
  OR2_X1 U1097 ( .A1(n138), .A2(n194), .ZN(n71) );
  OR2_X1 U1098 ( .A1(n154), .A2(n172), .ZN(n72) );
  OR2_X1 U1099 ( .A1(n138), .A2(n193), .ZN(n73) );
  OR2_X1 U1100 ( .A1(n138), .A2(n192), .ZN(n74) );
  OR2_X1 U1101 ( .A1(n136), .A2(n172), .ZN(n75) );
  OR2_X1 U1102 ( .A1(n138), .A2(n199), .ZN(n76) );
  OR2_X1 U1103 ( .A1(n138), .A2(n188), .ZN(n77) );
  OR2_X1 U1104 ( .A1(n153), .A2(n172), .ZN(n78) );
  OR2_X1 U1105 ( .A1(n168), .A2(n172), .ZN(n79) );
  OR2_X1 U1106 ( .A1(n167), .A2(n172), .ZN(n80) );
  OR2_X1 U1107 ( .A1(n152), .A2(n172), .ZN(n81) );
  OR2_X1 U1108 ( .A1(n138), .A2(n177), .ZN(n82) );
  OR2_X1 U1109 ( .A1(n138), .A2(n191), .ZN(n83) );
  OR2_X1 U1110 ( .A1(n166), .A2(n172), .ZN(n84) );
  OR2_X1 U1111 ( .A1(n138), .A2(n175), .ZN(n85) );
  OR2_X1 U1112 ( .A1(n138), .A2(n174), .ZN(n86) );
  OR2_X1 U1113 ( .A1(n165), .A2(n172), .ZN(n87) );
  OR2_X1 U1114 ( .A1(n164), .A2(n172), .ZN(n88) );
  OR2_X1 U1115 ( .A1(n138), .A2(n173), .ZN(n89) );
  OR2_X1 U1116 ( .A1(n163), .A2(n172), .ZN(n90) );
  OR2_X1 U1117 ( .A1(n138), .A2(n171), .ZN(n91) );
  OR2_X1 U1118 ( .A1(n138), .A2(n170), .ZN(n92) );
  OR2_X1 U1119 ( .A1(n162), .A2(n172), .ZN(n93) );
  OR2_X1 U1120 ( .A1(n161), .A2(n172), .ZN(n94) );
  OR2_X1 U1121 ( .A1(n138), .A2(n169), .ZN(n95) );
  OR2_X1 U1122 ( .A1(n160), .A2(n172), .ZN(n96) );
  OR2_X1 U1123 ( .A1(n137), .A2(n138), .ZN(n97) );
  OR2_X1 U1124 ( .A1(n138), .A2(n198), .ZN(n98) );
  INV_X2 U1125 ( .A(n83), .ZN(n99) );
  INV_X2 U1126 ( .A(n81), .ZN(n100) );
  INV_X2 U1127 ( .A(n78), .ZN(n101) );
  INV_X2 U1128 ( .A(n74), .ZN(n102) );
  INV_X2 U1129 ( .A(n73), .ZN(n103) );
  INV_X2 U1130 ( .A(n72), .ZN(n104) );
  INV_X2 U1131 ( .A(n71), .ZN(n105) );
  INV_X2 U1132 ( .A(n70), .ZN(n106) );
  INV_X2 U1133 ( .A(n69), .ZN(n107) );
  INV_X2 U1134 ( .A(n68), .ZN(n108) );
  INV_X2 U1135 ( .A(n67), .ZN(n109) );
  INV_X2 U1136 ( .A(n66), .ZN(n110) );
  INV_X2 U1137 ( .A(n64), .ZN(n111) );
  INV_X2 U1138 ( .A(n65), .ZN(n112) );
  INV_X4 U1139 ( .A(n98), .ZN(n113) );
  INV_X2 U1140 ( .A(n63), .ZN(n114) );
  INV_X4 U1141 ( .A(n96), .ZN(n115) );
  INV_X4 U1142 ( .A(n97), .ZN(n116) );
  INV_X4 U1143 ( .A(n94), .ZN(n117) );
  INV_X4 U1144 ( .A(n95), .ZN(n118) );
  INV_X4 U1145 ( .A(n92), .ZN(n119) );
  INV_X4 U1146 ( .A(n93), .ZN(n120) );
  INV_X4 U1147 ( .A(n90), .ZN(n121) );
  INV_X4 U1148 ( .A(n91), .ZN(n122) );
  INV_X4 U1149 ( .A(n88), .ZN(n123) );
  INV_X4 U1150 ( .A(n89), .ZN(n124) );
  INV_X4 U1151 ( .A(n86), .ZN(n125) );
  INV_X4 U1152 ( .A(n87), .ZN(n126) );
  INV_X4 U1153 ( .A(n84), .ZN(n127) );
  INV_X4 U1154 ( .A(n85), .ZN(n128) );
  INV_X4 U1155 ( .A(n80), .ZN(n129) );
  INV_X4 U1156 ( .A(n82), .ZN(n130) );
  INV_X4 U1157 ( .A(n77), .ZN(n131) );
  INV_X4 U1158 ( .A(n79), .ZN(n132) );
  INV_X4 U1159 ( .A(n75), .ZN(n133) );
  INV_X4 U1160 ( .A(n76), .ZN(n134) );
  NOR2_X2 U1161 ( .A1(n143), .A2(n172), .ZN(shiftedA_37__63_) );
  NOR2_X4 U1162 ( .A1(n149), .A2(n172), .ZN(shiftedA_43__63_) );
  NOR2_X2 U1163 ( .A1(n138), .A2(n181), .ZN(shiftedA_26__63_) );
  NOR2_X2 U1164 ( .A1(n144), .A2(n172), .ZN(shiftedA_38__63_) );
  NOR2_X2 U1165 ( .A1(n138), .A2(n184), .ZN(shiftedA_23__63_) );
  NOR2_X4 U1166 ( .A1(n147), .A2(n172), .ZN(shiftedA_41__63_) );
  NOR2_X4 U1167 ( .A1(n138), .A2(n187), .ZN(shiftedA_20__63_) );
  NOR2_X4 U1168 ( .A1(n150), .A2(n172), .ZN(shiftedA_44__63_) );
  NOR2_X2 U1169 ( .A1(n138), .A2(n183), .ZN(shiftedA_24__63_) );
  NOR2_X2 U1170 ( .A1(n145), .A2(n172), .ZN(shiftedA_39__63_) );
  NOR2_X4 U1171 ( .A1(n138), .A2(n185), .ZN(shiftedA_22__63_) );
  NOR2_X4 U1172 ( .A1(n148), .A2(n172), .ZN(shiftedA_42__63_) );
  NOR2_X4 U1173 ( .A1(n138), .A2(n189), .ZN(shiftedA_19__63_) );
  NOR2_X4 U1174 ( .A1(n151), .A2(n172), .ZN(shiftedA_45__63_) );
  NOR2_X2 U1175 ( .A1(n138), .A2(n182), .ZN(shiftedA_25__63_) );
  INV_X2 U1176 ( .A(b[30]), .ZN(n176) );
  INV_X2 U1177 ( .A(b[29]), .ZN(n178) );
  INV_X2 U1178 ( .A(b[28]), .ZN(n179) );
  INV_X2 U1179 ( .A(b[27]), .ZN(n180) );
  INV_X2 U1180 ( .A(b[26]), .ZN(n181) );
  INV_X2 U1181 ( .A(b[25]), .ZN(n182) );
  INV_X2 U1182 ( .A(b[24]), .ZN(n183) );
  INV_X2 U1183 ( .A(b[23]), .ZN(n184) );
  INV_X2 U1184 ( .A(b[22]), .ZN(n185) );
  INV_X2 U1185 ( .A(b[21]), .ZN(n186) );
  INV_X2 U1186 ( .A(b[20]), .ZN(n187) );
  INV_X2 U1187 ( .A(b[19]), .ZN(n189) );
  INV_X2 U1188 ( .A(b[18]), .ZN(n190) );
  INV_X2 U1189 ( .A(b[17]), .ZN(n191) );
  INV_X2 U1190 ( .A(b[16]), .ZN(n192) );
  INV_X2 U1191 ( .A(b[15]), .ZN(n193) );
  INV_X2 U1192 ( .A(b[14]), .ZN(n194) );
  INV_X2 U1193 ( .A(b[13]), .ZN(n195) );
  INV_X2 U1194 ( .A(b[12]), .ZN(n196) );
  INV_X2 U1195 ( .A(b[11]), .ZN(n197) );
  INV_X2 U1196 ( .A(b[10]), .ZN(n198) );
  INV_X2 U1197 ( .A(b[8]), .ZN(n169) );
  INV_X2 U1198 ( .A(b[7]), .ZN(n170) );
  INV_X2 U1199 ( .A(b[6]), .ZN(n171) );
  INV_X2 U1200 ( .A(b[5]), .ZN(n173) );
  INV_X2 U1201 ( .A(b[4]), .ZN(n174) );
  INV_X2 U1202 ( .A(b[3]), .ZN(n175) );
  INV_X2 U1203 ( .A(b[2]), .ZN(n177) );
  INV_X2 U1204 ( .A(b[1]), .ZN(n188) );
  INV_X2 U1205 ( .A(b[0]), .ZN(n199) );
  INV_X2 U1206 ( .A(b[31]), .ZN(n172) );
  NOR2_X2 U1207 ( .A1(n146), .A2(n172), .ZN(shiftedA_40__63_) );
  INV_X2 U1208 ( .A(a[30]), .ZN(n139) );
  INV_X2 U1209 ( .A(a[29]), .ZN(n140) );
  INV_X2 U1210 ( .A(a[28]), .ZN(n141) );
  INV_X2 U1211 ( .A(a[27]), .ZN(n142) );
  INV_X2 U1212 ( .A(a[26]), .ZN(n143) );
  INV_X2 U1213 ( .A(a[25]), .ZN(n144) );
  INV_X2 U1214 ( .A(a[24]), .ZN(n145) );
  INV_X2 U1215 ( .A(a[23]), .ZN(n146) );
  INV_X2 U1216 ( .A(a[22]), .ZN(n147) );
  INV_X2 U1217 ( .A(a[21]), .ZN(n148) );
  INV_X2 U1218 ( .A(a[20]), .ZN(n149) );
  INV_X2 U1219 ( .A(a[19]), .ZN(n150) );
  INV_X2 U1220 ( .A(a[18]), .ZN(n151) );
  INV_X2 U1221 ( .A(a[17]), .ZN(n152) );
  INV_X2 U1222 ( .A(a[16]), .ZN(n153) );
  INV_X2 U1223 ( .A(a[15]), .ZN(n154) );
  INV_X2 U1224 ( .A(a[14]), .ZN(n155) );
  INV_X2 U1225 ( .A(a[13]), .ZN(n156) );
  INV_X2 U1226 ( .A(a[11]), .ZN(n158) );
  INV_X2 U1227 ( .A(a[12]), .ZN(n157) );
  INV_X2 U1228 ( .A(a[10]), .ZN(n159) );
  INV_X2 U1229 ( .A(b[9]), .ZN(n137) );
  INV_X2 U1230 ( .A(a[9]), .ZN(n160) );
  INV_X2 U1231 ( .A(a[8]), .ZN(n161) );
  INV_X2 U1232 ( .A(a[7]), .ZN(n162) );
  INV_X2 U1233 ( .A(a[6]), .ZN(n163) );
  INV_X2 U1234 ( .A(a[5]), .ZN(n164) );
  INV_X2 U1235 ( .A(a[4]), .ZN(n165) );
  INV_X2 U1236 ( .A(a[3]), .ZN(n166) );
  INV_X2 U1237 ( .A(a[2]), .ZN(n167) );
  INV_X2 U1238 ( .A(a[1]), .ZN(n168) );
  INV_X2 U1239 ( .A(a[31]), .ZN(n138) );
  INV_X2 U1240 ( .A(a[0]), .ZN(n136) );
  NOR2_X4 U1241 ( .A1(n138), .A2(n186), .ZN(shiftedA_21__63_) );
  NOR2_X4 U1242 ( .A1(n138), .A2(n190), .ZN(shiftedA_18__63_) );
  NOR2_X1 U1244 ( .A1(n136), .A2(n137), .ZN(shiftedA_9__9_) );
  NOR2_X1 U1245 ( .A1(n137), .A2(n139), .ZN(shiftedA_9__39_) );
  NOR2_X1 U1246 ( .A1(n137), .A2(n140), .ZN(shiftedA_9__38_) );
  NOR2_X1 U1247 ( .A1(n137), .A2(n141), .ZN(shiftedA_9__37_) );
  NOR2_X1 U1248 ( .A1(n137), .A2(n142), .ZN(shiftedA_9__36_) );
  NOR2_X1 U1249 ( .A1(n137), .A2(n143), .ZN(shiftedA_9__35_) );
  NOR2_X1 U1250 ( .A1(n137), .A2(n144), .ZN(shiftedA_9__34_) );
  NOR2_X1 U1251 ( .A1(n137), .A2(n145), .ZN(shiftedA_9__33_) );
  NOR2_X1 U1252 ( .A1(n137), .A2(n146), .ZN(shiftedA_9__32_) );
  NOR2_X1 U1253 ( .A1(n137), .A2(n147), .ZN(shiftedA_9__31_) );
  NOR2_X1 U1254 ( .A1(n137), .A2(n148), .ZN(shiftedA_9__30_) );
  NOR2_X1 U1255 ( .A1(n137), .A2(n149), .ZN(shiftedA_9__29_) );
  NOR2_X1 U1256 ( .A1(n137), .A2(n150), .ZN(shiftedA_9__28_) );
  NOR2_X1 U1257 ( .A1(n137), .A2(n151), .ZN(shiftedA_9__27_) );
  NOR2_X1 U1258 ( .A1(n137), .A2(n152), .ZN(shiftedA_9__26_) );
  NOR2_X1 U1259 ( .A1(n137), .A2(n153), .ZN(shiftedA_9__25_) );
  NOR2_X1 U1260 ( .A1(n137), .A2(n154), .ZN(shiftedA_9__24_) );
  NOR2_X1 U1261 ( .A1(n137), .A2(n155), .ZN(shiftedA_9__23_) );
  NOR2_X1 U1262 ( .A1(n137), .A2(n156), .ZN(shiftedA_9__22_) );
  NOR2_X1 U1263 ( .A1(n137), .A2(n157), .ZN(shiftedA_9__21_) );
  NOR2_X1 U1264 ( .A1(n137), .A2(n158), .ZN(shiftedA_9__20_) );
  NOR2_X1 U1265 ( .A1(n137), .A2(n159), .ZN(shiftedA_9__19_) );
  NOR2_X1 U1266 ( .A1(n137), .A2(n160), .ZN(shiftedA_9__18_) );
  NOR2_X1 U1267 ( .A1(n137), .A2(n161), .ZN(shiftedA_9__17_) );
  NOR2_X1 U1268 ( .A1(n137), .A2(n162), .ZN(shiftedA_9__16_) );
  NOR2_X1 U1269 ( .A1(n137), .A2(n163), .ZN(shiftedA_9__15_) );
  NOR2_X1 U1270 ( .A1(n137), .A2(n164), .ZN(shiftedA_9__14_) );
  NOR2_X1 U1271 ( .A1(n137), .A2(n165), .ZN(shiftedA_9__13_) );
  NOR2_X1 U1272 ( .A1(n137), .A2(n166), .ZN(shiftedA_9__12_) );
  NOR2_X1 U1273 ( .A1(n137), .A2(n167), .ZN(shiftedA_9__11_) );
  NOR2_X1 U1274 ( .A1(n137), .A2(n168), .ZN(shiftedA_9__10_) );
  NOR2_X1 U1275 ( .A1(n168), .A2(n169), .ZN(shiftedA_8__9_) );
  NOR2_X1 U1276 ( .A1(n136), .A2(n169), .ZN(shiftedA_8__8_) );
  NOR2_X1 U1277 ( .A1(n139), .A2(n169), .ZN(shiftedA_8__38_) );
  NOR2_X1 U1278 ( .A1(n140), .A2(n169), .ZN(shiftedA_8__37_) );
  NOR2_X1 U1279 ( .A1(n141), .A2(n169), .ZN(shiftedA_8__36_) );
  NOR2_X1 U1280 ( .A1(n142), .A2(n169), .ZN(shiftedA_8__35_) );
  NOR2_X1 U1281 ( .A1(n143), .A2(n169), .ZN(shiftedA_8__34_) );
  NOR2_X1 U1282 ( .A1(n144), .A2(n169), .ZN(shiftedA_8__33_) );
  NOR2_X1 U1283 ( .A1(n145), .A2(n169), .ZN(shiftedA_8__32_) );
  NOR2_X1 U1284 ( .A1(n146), .A2(n169), .ZN(shiftedA_8__31_) );
  NOR2_X1 U1285 ( .A1(n147), .A2(n169), .ZN(shiftedA_8__30_) );
  NOR2_X1 U1286 ( .A1(n148), .A2(n169), .ZN(shiftedA_8__29_) );
  NOR2_X1 U1287 ( .A1(n149), .A2(n169), .ZN(shiftedA_8__28_) );
  NOR2_X1 U1288 ( .A1(n150), .A2(n169), .ZN(shiftedA_8__27_) );
  NOR2_X1 U1289 ( .A1(n151), .A2(n169), .ZN(shiftedA_8__26_) );
  NOR2_X1 U1290 ( .A1(n152), .A2(n169), .ZN(shiftedA_8__25_) );
  NOR2_X1 U1291 ( .A1(n153), .A2(n169), .ZN(shiftedA_8__24_) );
  NOR2_X1 U1292 ( .A1(n154), .A2(n169), .ZN(shiftedA_8__23_) );
  NOR2_X1 U1293 ( .A1(n155), .A2(n169), .ZN(shiftedA_8__22_) );
  NOR2_X1 U1294 ( .A1(n156), .A2(n169), .ZN(shiftedA_8__21_) );
  NOR2_X1 U1295 ( .A1(n157), .A2(n169), .ZN(shiftedA_8__20_) );
  NOR2_X1 U1296 ( .A1(n158), .A2(n169), .ZN(shiftedA_8__19_) );
  NOR2_X1 U1297 ( .A1(n159), .A2(n169), .ZN(shiftedA_8__18_) );
  NOR2_X1 U1298 ( .A1(n160), .A2(n169), .ZN(shiftedA_8__17_) );
  NOR2_X1 U1299 ( .A1(n161), .A2(n169), .ZN(shiftedA_8__16_) );
  NOR2_X1 U1300 ( .A1(n162), .A2(n169), .ZN(shiftedA_8__15_) );
  NOR2_X1 U1301 ( .A1(n163), .A2(n169), .ZN(shiftedA_8__14_) );
  NOR2_X1 U1302 ( .A1(n164), .A2(n169), .ZN(shiftedA_8__13_) );
  NOR2_X1 U1303 ( .A1(n165), .A2(n169), .ZN(shiftedA_8__12_) );
  NOR2_X1 U1304 ( .A1(n166), .A2(n169), .ZN(shiftedA_8__11_) );
  NOR2_X1 U1305 ( .A1(n167), .A2(n169), .ZN(shiftedA_8__10_) );
  NOR2_X1 U1306 ( .A1(n167), .A2(n170), .ZN(shiftedA_7__9_) );
  NOR2_X1 U1307 ( .A1(n168), .A2(n170), .ZN(shiftedA_7__8_) );
  NOR2_X1 U1308 ( .A1(n136), .A2(n170), .ZN(shiftedA_7__7_) );
  NOR2_X1 U1309 ( .A1(n139), .A2(n170), .ZN(shiftedA_7__37_) );
  NOR2_X1 U1310 ( .A1(n140), .A2(n170), .ZN(shiftedA_7__36_) );
  NOR2_X1 U1311 ( .A1(n141), .A2(n170), .ZN(shiftedA_7__35_) );
  NOR2_X1 U1312 ( .A1(n142), .A2(n170), .ZN(shiftedA_7__34_) );
  NOR2_X1 U1313 ( .A1(n143), .A2(n170), .ZN(shiftedA_7__33_) );
  NOR2_X1 U1314 ( .A1(n144), .A2(n170), .ZN(shiftedA_7__32_) );
  NOR2_X1 U1315 ( .A1(n145), .A2(n170), .ZN(shiftedA_7__31_) );
  NOR2_X1 U1316 ( .A1(n146), .A2(n170), .ZN(shiftedA_7__30_) );
  NOR2_X1 U1317 ( .A1(n147), .A2(n170), .ZN(shiftedA_7__29_) );
  NOR2_X1 U1318 ( .A1(n148), .A2(n170), .ZN(shiftedA_7__28_) );
  NOR2_X1 U1319 ( .A1(n149), .A2(n170), .ZN(shiftedA_7__27_) );
  NOR2_X1 U1320 ( .A1(n150), .A2(n170), .ZN(shiftedA_7__26_) );
  NOR2_X1 U1321 ( .A1(n151), .A2(n170), .ZN(shiftedA_7__25_) );
  NOR2_X1 U1322 ( .A1(n152), .A2(n170), .ZN(shiftedA_7__24_) );
  NOR2_X1 U1323 ( .A1(n153), .A2(n170), .ZN(shiftedA_7__23_) );
  NOR2_X1 U1324 ( .A1(n154), .A2(n170), .ZN(shiftedA_7__22_) );
  NOR2_X1 U1325 ( .A1(n155), .A2(n170), .ZN(shiftedA_7__21_) );
  NOR2_X1 U1326 ( .A1(n156), .A2(n170), .ZN(shiftedA_7__20_) );
  NOR2_X1 U1327 ( .A1(n157), .A2(n170), .ZN(shiftedA_7__19_) );
  NOR2_X1 U1328 ( .A1(n158), .A2(n170), .ZN(shiftedA_7__18_) );
  NOR2_X1 U1329 ( .A1(n159), .A2(n170), .ZN(shiftedA_7__17_) );
  NOR2_X1 U1330 ( .A1(n160), .A2(n170), .ZN(shiftedA_7__16_) );
  NOR2_X1 U1331 ( .A1(n161), .A2(n170), .ZN(shiftedA_7__15_) );
  NOR2_X1 U1332 ( .A1(n162), .A2(n170), .ZN(shiftedA_7__14_) );
  NOR2_X1 U1333 ( .A1(n163), .A2(n170), .ZN(shiftedA_7__13_) );
  NOR2_X1 U1334 ( .A1(n164), .A2(n170), .ZN(shiftedA_7__12_) );
  NOR2_X1 U1335 ( .A1(n165), .A2(n170), .ZN(shiftedA_7__11_) );
  NOR2_X1 U1336 ( .A1(n166), .A2(n170), .ZN(shiftedA_7__10_) );
  NOR2_X1 U1337 ( .A1(n166), .A2(n171), .ZN(shiftedA_6__9_) );
  NOR2_X1 U1338 ( .A1(n167), .A2(n171), .ZN(shiftedA_6__8_) );
  NOR2_X1 U1339 ( .A1(n168), .A2(n171), .ZN(shiftedA_6__7_) );
  NOR2_X1 U1340 ( .A1(n136), .A2(n171), .ZN(shiftedA_6__6_) );
  NOR2_X1 U1341 ( .A1(n139), .A2(n171), .ZN(shiftedA_6__36_) );
  NOR2_X1 U1342 ( .A1(n140), .A2(n171), .ZN(shiftedA_6__35_) );
  NOR2_X1 U1343 ( .A1(n141), .A2(n171), .ZN(shiftedA_6__34_) );
  NOR2_X1 U1344 ( .A1(n142), .A2(n171), .ZN(shiftedA_6__33_) );
  NOR2_X1 U1345 ( .A1(n143), .A2(n171), .ZN(shiftedA_6__32_) );
  NOR2_X1 U1346 ( .A1(n144), .A2(n171), .ZN(shiftedA_6__31_) );
  NOR2_X1 U1347 ( .A1(n145), .A2(n171), .ZN(shiftedA_6__30_) );
  NOR2_X1 U1348 ( .A1(n146), .A2(n171), .ZN(shiftedA_6__29_) );
  NOR2_X1 U1349 ( .A1(n147), .A2(n171), .ZN(shiftedA_6__28_) );
  NOR2_X1 U1350 ( .A1(n148), .A2(n171), .ZN(shiftedA_6__27_) );
  NOR2_X1 U1351 ( .A1(n149), .A2(n171), .ZN(shiftedA_6__26_) );
  NOR2_X1 U1352 ( .A1(n150), .A2(n171), .ZN(shiftedA_6__25_) );
  NOR2_X1 U1353 ( .A1(n151), .A2(n171), .ZN(shiftedA_6__24_) );
  NOR2_X1 U1354 ( .A1(n152), .A2(n171), .ZN(shiftedA_6__23_) );
  NOR2_X1 U1355 ( .A1(n153), .A2(n171), .ZN(shiftedA_6__22_) );
  NOR2_X1 U1356 ( .A1(n154), .A2(n171), .ZN(shiftedA_6__21_) );
  NOR2_X1 U1357 ( .A1(n155), .A2(n171), .ZN(shiftedA_6__20_) );
  NOR2_X1 U1358 ( .A1(n156), .A2(n171), .ZN(shiftedA_6__19_) );
  NOR2_X1 U1359 ( .A1(n157), .A2(n171), .ZN(shiftedA_6__18_) );
  NOR2_X1 U1360 ( .A1(n158), .A2(n171), .ZN(shiftedA_6__17_) );
  NOR2_X1 U1361 ( .A1(n159), .A2(n171), .ZN(shiftedA_6__16_) );
  NOR2_X1 U1362 ( .A1(n160), .A2(n171), .ZN(shiftedA_6__15_) );
  NOR2_X1 U1363 ( .A1(n161), .A2(n171), .ZN(shiftedA_6__14_) );
  NOR2_X1 U1364 ( .A1(n162), .A2(n171), .ZN(shiftedA_6__13_) );
  NOR2_X1 U1365 ( .A1(n163), .A2(n171), .ZN(shiftedA_6__12_) );
  NOR2_X1 U1366 ( .A1(n164), .A2(n171), .ZN(shiftedA_6__11_) );
  NOR2_X1 U1367 ( .A1(n165), .A2(n171), .ZN(shiftedA_6__10_) );
  NOR2_X1 U1368 ( .A1(n165), .A2(n173), .ZN(shiftedA_5__9_) );
  NOR2_X1 U1369 ( .A1(n166), .A2(n173), .ZN(shiftedA_5__8_) );
  NOR2_X1 U1370 ( .A1(n167), .A2(n173), .ZN(shiftedA_5__7_) );
  NOR2_X1 U1371 ( .A1(n168), .A2(n173), .ZN(shiftedA_5__6_) );
  NOR2_X1 U1372 ( .A1(n136), .A2(n173), .ZN(shiftedA_5__5_) );
  NOR2_X1 U1373 ( .A1(n139), .A2(n173), .ZN(shiftedA_5__35_) );
  NOR2_X1 U1374 ( .A1(n140), .A2(n173), .ZN(shiftedA_5__34_) );
  NOR2_X1 U1375 ( .A1(n141), .A2(n173), .ZN(shiftedA_5__33_) );
  NOR2_X1 U1376 ( .A1(n142), .A2(n173), .ZN(shiftedA_5__32_) );
  NOR2_X1 U1377 ( .A1(n143), .A2(n173), .ZN(shiftedA_5__31_) );
  NOR2_X1 U1378 ( .A1(n144), .A2(n173), .ZN(shiftedA_5__30_) );
  NOR2_X1 U1379 ( .A1(n145), .A2(n173), .ZN(shiftedA_5__29_) );
  NOR2_X1 U1380 ( .A1(n146), .A2(n173), .ZN(shiftedA_5__28_) );
  NOR2_X1 U1381 ( .A1(n147), .A2(n173), .ZN(shiftedA_5__27_) );
  NOR2_X1 U1382 ( .A1(n148), .A2(n173), .ZN(shiftedA_5__26_) );
  NOR2_X1 U1383 ( .A1(n149), .A2(n173), .ZN(shiftedA_5__25_) );
  NOR2_X1 U1384 ( .A1(n150), .A2(n173), .ZN(shiftedA_5__24_) );
  NOR2_X1 U1385 ( .A1(n151), .A2(n173), .ZN(shiftedA_5__23_) );
  NOR2_X1 U1386 ( .A1(n152), .A2(n173), .ZN(shiftedA_5__22_) );
  NOR2_X1 U1387 ( .A1(n153), .A2(n173), .ZN(shiftedA_5__21_) );
  NOR2_X1 U1388 ( .A1(n154), .A2(n173), .ZN(shiftedA_5__20_) );
  NOR2_X1 U1389 ( .A1(n155), .A2(n173), .ZN(shiftedA_5__19_) );
  NOR2_X1 U1390 ( .A1(n156), .A2(n173), .ZN(shiftedA_5__18_) );
  NOR2_X1 U1391 ( .A1(n157), .A2(n173), .ZN(shiftedA_5__17_) );
  NOR2_X1 U1392 ( .A1(n158), .A2(n173), .ZN(shiftedA_5__16_) );
  NOR2_X1 U1393 ( .A1(n159), .A2(n173), .ZN(shiftedA_5__15_) );
  NOR2_X1 U1394 ( .A1(n160), .A2(n173), .ZN(shiftedA_5__14_) );
  NOR2_X1 U1395 ( .A1(n161), .A2(n173), .ZN(shiftedA_5__13_) );
  NOR2_X1 U1396 ( .A1(n162), .A2(n173), .ZN(shiftedA_5__12_) );
  NOR2_X1 U1397 ( .A1(n163), .A2(n173), .ZN(shiftedA_5__11_) );
  NOR2_X1 U1398 ( .A1(n164), .A2(n173), .ZN(shiftedA_5__10_) );
  NOR2_X1 U1399 ( .A1(n164), .A2(n174), .ZN(shiftedA_4__9_) );
  NOR2_X1 U1400 ( .A1(n165), .A2(n174), .ZN(shiftedA_4__8_) );
  NOR2_X1 U1401 ( .A1(n166), .A2(n174), .ZN(shiftedA_4__7_) );
  NOR2_X1 U1402 ( .A1(n167), .A2(n174), .ZN(shiftedA_4__6_) );
  NOR2_X1 U1403 ( .A1(n168), .A2(n174), .ZN(shiftedA_4__5_) );
  NOR2_X1 U1404 ( .A1(n136), .A2(n174), .ZN(shiftedA_4__4_) );
  NOR2_X1 U1405 ( .A1(n139), .A2(n174), .ZN(shiftedA_4__34_) );
  NOR2_X1 U1406 ( .A1(n140), .A2(n174), .ZN(shiftedA_4__33_) );
  NOR2_X1 U1407 ( .A1(n141), .A2(n174), .ZN(shiftedA_4__32_) );
  NOR2_X1 U1408 ( .A1(n142), .A2(n174), .ZN(shiftedA_4__31_) );
  NOR2_X1 U1409 ( .A1(n143), .A2(n174), .ZN(shiftedA_4__30_) );
  NOR2_X1 U1410 ( .A1(n144), .A2(n174), .ZN(shiftedA_4__29_) );
  NOR2_X1 U1411 ( .A1(n145), .A2(n174), .ZN(shiftedA_4__28_) );
  NOR2_X1 U1412 ( .A1(n146), .A2(n174), .ZN(shiftedA_4__27_) );
  NOR2_X1 U1413 ( .A1(n147), .A2(n174), .ZN(shiftedA_4__26_) );
  NOR2_X1 U1414 ( .A1(n148), .A2(n174), .ZN(shiftedA_4__25_) );
  NOR2_X1 U1415 ( .A1(n149), .A2(n174), .ZN(shiftedA_4__24_) );
  NOR2_X1 U1416 ( .A1(n150), .A2(n174), .ZN(shiftedA_4__23_) );
  NOR2_X1 U1417 ( .A1(n151), .A2(n174), .ZN(shiftedA_4__22_) );
  NOR2_X1 U1418 ( .A1(n152), .A2(n174), .ZN(shiftedA_4__21_) );
  NOR2_X1 U1419 ( .A1(n153), .A2(n174), .ZN(shiftedA_4__20_) );
  NOR2_X1 U1420 ( .A1(n154), .A2(n174), .ZN(shiftedA_4__19_) );
  NOR2_X1 U1421 ( .A1(n155), .A2(n174), .ZN(shiftedA_4__18_) );
  NOR2_X1 U1422 ( .A1(n156), .A2(n174), .ZN(shiftedA_4__17_) );
  NOR2_X1 U1423 ( .A1(n157), .A2(n174), .ZN(shiftedA_4__16_) );
  NOR2_X1 U1424 ( .A1(n158), .A2(n174), .ZN(shiftedA_4__15_) );
  NOR2_X1 U1425 ( .A1(n159), .A2(n174), .ZN(shiftedA_4__14_) );
  NOR2_X1 U1426 ( .A1(n160), .A2(n174), .ZN(shiftedA_4__13_) );
  NOR2_X1 U1427 ( .A1(n161), .A2(n174), .ZN(shiftedA_4__12_) );
  NOR2_X1 U1428 ( .A1(n162), .A2(n174), .ZN(shiftedA_4__11_) );
  NOR2_X1 U1429 ( .A1(n163), .A2(n174), .ZN(shiftedA_4__10_) );
  NOR2_X1 U1430 ( .A1(n163), .A2(n175), .ZN(shiftedA_3__9_) );
  NOR2_X1 U1431 ( .A1(n164), .A2(n175), .ZN(shiftedA_3__8_) );
  NOR2_X1 U1432 ( .A1(n165), .A2(n175), .ZN(shiftedA_3__7_) );
  NOR2_X1 U1433 ( .A1(n166), .A2(n175), .ZN(shiftedA_3__6_) );
  NOR2_X1 U1434 ( .A1(n167), .A2(n175), .ZN(shiftedA_3__5_) );
  NOR2_X1 U1435 ( .A1(n168), .A2(n175), .ZN(shiftedA_3__4_) );
  NOR2_X1 U1436 ( .A1(n136), .A2(n175), .ZN(shiftedA_3__3_) );
  NOR2_X1 U1437 ( .A1(n139), .A2(n175), .ZN(shiftedA_3__33_) );
  NOR2_X1 U1438 ( .A1(n140), .A2(n175), .ZN(shiftedA_3__32_) );
  NOR2_X1 U1439 ( .A1(n141), .A2(n175), .ZN(shiftedA_3__31_) );
  NOR2_X1 U1440 ( .A1(n142), .A2(n175), .ZN(shiftedA_3__30_) );
  NOR2_X1 U1441 ( .A1(n143), .A2(n175), .ZN(shiftedA_3__29_) );
  NOR2_X1 U1442 ( .A1(n144), .A2(n175), .ZN(shiftedA_3__28_) );
  NOR2_X1 U1443 ( .A1(n145), .A2(n175), .ZN(shiftedA_3__27_) );
  NOR2_X1 U1444 ( .A1(n146), .A2(n175), .ZN(shiftedA_3__26_) );
  NOR2_X1 U1445 ( .A1(n147), .A2(n175), .ZN(shiftedA_3__25_) );
  NOR2_X1 U1446 ( .A1(n148), .A2(n175), .ZN(shiftedA_3__24_) );
  NOR2_X1 U1447 ( .A1(n149), .A2(n175), .ZN(shiftedA_3__23_) );
  NOR2_X1 U1448 ( .A1(n150), .A2(n175), .ZN(shiftedA_3__22_) );
  NOR2_X1 U1449 ( .A1(n151), .A2(n175), .ZN(shiftedA_3__21_) );
  NOR2_X1 U1450 ( .A1(n152), .A2(n175), .ZN(shiftedA_3__20_) );
  NOR2_X1 U1451 ( .A1(n153), .A2(n175), .ZN(shiftedA_3__19_) );
  NOR2_X1 U1452 ( .A1(n154), .A2(n175), .ZN(shiftedA_3__18_) );
  NOR2_X1 U1453 ( .A1(n155), .A2(n175), .ZN(shiftedA_3__17_) );
  NOR2_X1 U1454 ( .A1(n156), .A2(n175), .ZN(shiftedA_3__16_) );
  NOR2_X1 U1455 ( .A1(n157), .A2(n175), .ZN(shiftedA_3__15_) );
  NOR2_X1 U1456 ( .A1(n158), .A2(n175), .ZN(shiftedA_3__14_) );
  NOR2_X1 U1457 ( .A1(n159), .A2(n175), .ZN(shiftedA_3__13_) );
  NOR2_X1 U1458 ( .A1(n160), .A2(n175), .ZN(shiftedA_3__12_) );
  NOR2_X1 U1459 ( .A1(n161), .A2(n175), .ZN(shiftedA_3__11_) );
  NOR2_X1 U1460 ( .A1(n162), .A2(n175), .ZN(shiftedA_3__10_) );
  NOR2_X1 U1461 ( .A1(n142), .A2(n172), .ZN(shiftedA_36__63_) );
  NOR2_X1 U1462 ( .A1(n141), .A2(n172), .ZN(shiftedA_35__63_) );
  NOR2_X1 U1463 ( .A1(n140), .A2(n172), .ZN(shiftedA_34__63_) );
  NOR2_X1 U1464 ( .A1(n139), .A2(n172), .ZN(shiftedA_33__63_) );
  NOR2_X1 U1465 ( .A1(n138), .A2(n172), .ZN(shiftedA_32__63_) );
  NOR2_X1 U1466 ( .A1(n138), .A2(n176), .ZN(shiftedA_30__63_) );
  NOR2_X1 U1467 ( .A1(n139), .A2(n176), .ZN(shiftedA_30__60_) );
  NOR2_X1 U1468 ( .A1(n140), .A2(n176), .ZN(shiftedA_30__59_) );
  NOR2_X1 U1469 ( .A1(n141), .A2(n176), .ZN(shiftedA_30__58_) );
  NOR2_X1 U1470 ( .A1(n142), .A2(n176), .ZN(shiftedA_30__57_) );
  NOR2_X1 U1471 ( .A1(n143), .A2(n176), .ZN(shiftedA_30__56_) );
  NOR2_X1 U1472 ( .A1(n144), .A2(n176), .ZN(shiftedA_30__55_) );
  NOR2_X1 U1473 ( .A1(n145), .A2(n176), .ZN(shiftedA_30__54_) );
  NOR2_X1 U1474 ( .A1(n146), .A2(n176), .ZN(shiftedA_30__53_) );
  NOR2_X1 U1475 ( .A1(n147), .A2(n176), .ZN(shiftedA_30__52_) );
  NOR2_X1 U1476 ( .A1(n148), .A2(n176), .ZN(shiftedA_30__51_) );
  NOR2_X1 U1477 ( .A1(n149), .A2(n176), .ZN(shiftedA_30__50_) );
  NOR2_X1 U1478 ( .A1(n150), .A2(n176), .ZN(shiftedA_30__49_) );
  NOR2_X1 U1479 ( .A1(n151), .A2(n176), .ZN(shiftedA_30__48_) );
  NOR2_X1 U1480 ( .A1(n152), .A2(n176), .ZN(shiftedA_30__47_) );
  NOR2_X1 U1481 ( .A1(n153), .A2(n176), .ZN(shiftedA_30__46_) );
  NOR2_X1 U1482 ( .A1(n154), .A2(n176), .ZN(shiftedA_30__45_) );
  NOR2_X1 U1483 ( .A1(n155), .A2(n176), .ZN(shiftedA_30__44_) );
  NOR2_X1 U1484 ( .A1(n156), .A2(n176), .ZN(shiftedA_30__43_) );
  NOR2_X1 U1485 ( .A1(n157), .A2(n176), .ZN(shiftedA_30__42_) );
  NOR2_X1 U1486 ( .A1(n158), .A2(n176), .ZN(shiftedA_30__41_) );
  NOR2_X1 U1487 ( .A1(n159), .A2(n176), .ZN(shiftedA_30__40_) );
  NOR2_X1 U1488 ( .A1(n160), .A2(n176), .ZN(shiftedA_30__39_) );
  NOR2_X1 U1489 ( .A1(n161), .A2(n176), .ZN(shiftedA_30__38_) );
  NOR2_X1 U1490 ( .A1(n162), .A2(n176), .ZN(shiftedA_30__37_) );
  NOR2_X1 U1491 ( .A1(n163), .A2(n176), .ZN(shiftedA_30__36_) );
  NOR2_X1 U1492 ( .A1(n164), .A2(n176), .ZN(shiftedA_30__35_) );
  NOR2_X1 U1493 ( .A1(n165), .A2(n176), .ZN(shiftedA_30__34_) );
  NOR2_X1 U1494 ( .A1(n166), .A2(n176), .ZN(shiftedA_30__33_) );
  NOR2_X1 U1495 ( .A1(n167), .A2(n176), .ZN(shiftedA_30__32_) );
  NOR2_X1 U1496 ( .A1(n168), .A2(n176), .ZN(shiftedA_30__31_) );
  NOR2_X1 U1497 ( .A1(n136), .A2(n176), .ZN(shiftedA_30__30_) );
  NOR2_X1 U1498 ( .A1(n162), .A2(n177), .ZN(shiftedA_2__9_) );
  NOR2_X1 U1499 ( .A1(n163), .A2(n177), .ZN(shiftedA_2__8_) );
  NOR2_X1 U1500 ( .A1(n164), .A2(n177), .ZN(shiftedA_2__7_) );
  NOR2_X1 U1501 ( .A1(n165), .A2(n177), .ZN(shiftedA_2__6_) );
  NOR2_X1 U1502 ( .A1(n166), .A2(n177), .ZN(shiftedA_2__5_) );
  NOR2_X1 U1503 ( .A1(n167), .A2(n177), .ZN(shiftedA_2__4_) );
  NOR2_X1 U1504 ( .A1(n168), .A2(n177), .ZN(shiftedA_2__3_) );
  NOR2_X1 U1505 ( .A1(n139), .A2(n177), .ZN(shiftedA_2__32_) );
  NOR2_X1 U1506 ( .A1(n140), .A2(n177), .ZN(shiftedA_2__31_) );
  NOR2_X1 U1507 ( .A1(n141), .A2(n177), .ZN(shiftedA_2__30_) );
  NOR2_X1 U1508 ( .A1(n136), .A2(n177), .ZN(shiftedA_2__2_) );
  NOR2_X1 U1509 ( .A1(n142), .A2(n177), .ZN(shiftedA_2__29_) );
  NOR2_X1 U1510 ( .A1(n143), .A2(n177), .ZN(shiftedA_2__28_) );
  NOR2_X1 U1511 ( .A1(n144), .A2(n177), .ZN(shiftedA_2__27_) );
  NOR2_X1 U1512 ( .A1(n145), .A2(n177), .ZN(shiftedA_2__26_) );
  NOR2_X1 U1513 ( .A1(n146), .A2(n177), .ZN(shiftedA_2__25_) );
  NOR2_X1 U1514 ( .A1(n147), .A2(n177), .ZN(shiftedA_2__24_) );
  NOR2_X1 U1515 ( .A1(n148), .A2(n177), .ZN(shiftedA_2__23_) );
  NOR2_X1 U1516 ( .A1(n149), .A2(n177), .ZN(shiftedA_2__22_) );
  NOR2_X1 U1517 ( .A1(n150), .A2(n177), .ZN(shiftedA_2__21_) );
  NOR2_X1 U1518 ( .A1(n151), .A2(n177), .ZN(shiftedA_2__20_) );
  NOR2_X1 U1519 ( .A1(n152), .A2(n177), .ZN(shiftedA_2__19_) );
  NOR2_X1 U1520 ( .A1(n153), .A2(n177), .ZN(shiftedA_2__18_) );
  NOR2_X1 U1521 ( .A1(n154), .A2(n177), .ZN(shiftedA_2__17_) );
  NOR2_X1 U1522 ( .A1(n155), .A2(n177), .ZN(shiftedA_2__16_) );
  NOR2_X1 U1523 ( .A1(n156), .A2(n177), .ZN(shiftedA_2__15_) );
  NOR2_X1 U1524 ( .A1(n157), .A2(n177), .ZN(shiftedA_2__14_) );
  NOR2_X1 U1525 ( .A1(n158), .A2(n177), .ZN(shiftedA_2__13_) );
  NOR2_X1 U1526 ( .A1(n159), .A2(n177), .ZN(shiftedA_2__12_) );
  NOR2_X1 U1527 ( .A1(n160), .A2(n177), .ZN(shiftedA_2__11_) );
  NOR2_X1 U1528 ( .A1(n161), .A2(n177), .ZN(shiftedA_2__10_) );
  NOR2_X1 U1529 ( .A1(n138), .A2(n178), .ZN(shiftedA_29__63_) );
  NOR2_X1 U1530 ( .A1(n139), .A2(n178), .ZN(shiftedA_29__59_) );
  NOR2_X1 U1531 ( .A1(n140), .A2(n178), .ZN(shiftedA_29__58_) );
  NOR2_X1 U1532 ( .A1(n141), .A2(n178), .ZN(shiftedA_29__57_) );
  NOR2_X1 U1533 ( .A1(n142), .A2(n178), .ZN(shiftedA_29__56_) );
  NOR2_X1 U1534 ( .A1(n143), .A2(n178), .ZN(shiftedA_29__55_) );
  NOR2_X1 U1535 ( .A1(n144), .A2(n178), .ZN(shiftedA_29__54_) );
  NOR2_X1 U1536 ( .A1(n145), .A2(n178), .ZN(shiftedA_29__53_) );
  NOR2_X1 U1537 ( .A1(n146), .A2(n178), .ZN(shiftedA_29__52_) );
  NOR2_X1 U1538 ( .A1(n147), .A2(n178), .ZN(shiftedA_29__51_) );
  NOR2_X1 U1539 ( .A1(n148), .A2(n178), .ZN(shiftedA_29__50_) );
  NOR2_X1 U1540 ( .A1(n149), .A2(n178), .ZN(shiftedA_29__49_) );
  NOR2_X1 U1541 ( .A1(n150), .A2(n178), .ZN(shiftedA_29__48_) );
  NOR2_X1 U1542 ( .A1(n151), .A2(n178), .ZN(shiftedA_29__47_) );
  NOR2_X1 U1543 ( .A1(n152), .A2(n178), .ZN(shiftedA_29__46_) );
  NOR2_X1 U1544 ( .A1(n153), .A2(n178), .ZN(shiftedA_29__45_) );
  NOR2_X1 U1545 ( .A1(n154), .A2(n178), .ZN(shiftedA_29__44_) );
  NOR2_X1 U1546 ( .A1(n155), .A2(n178), .ZN(shiftedA_29__43_) );
  NOR2_X1 U1547 ( .A1(n156), .A2(n178), .ZN(shiftedA_29__42_) );
  NOR2_X1 U1548 ( .A1(n157), .A2(n178), .ZN(shiftedA_29__41_) );
  NOR2_X1 U1549 ( .A1(n158), .A2(n178), .ZN(shiftedA_29__40_) );
  NOR2_X1 U1550 ( .A1(n159), .A2(n178), .ZN(shiftedA_29__39_) );
  NOR2_X1 U1551 ( .A1(n160), .A2(n178), .ZN(shiftedA_29__38_) );
  NOR2_X1 U1552 ( .A1(n161), .A2(n178), .ZN(shiftedA_29__37_) );
  NOR2_X1 U1553 ( .A1(n162), .A2(n178), .ZN(shiftedA_29__36_) );
  NOR2_X1 U1554 ( .A1(n163), .A2(n178), .ZN(shiftedA_29__35_) );
  NOR2_X1 U1555 ( .A1(n164), .A2(n178), .ZN(shiftedA_29__34_) );
  NOR2_X1 U1556 ( .A1(n165), .A2(n178), .ZN(shiftedA_29__33_) );
  NOR2_X1 U1557 ( .A1(n166), .A2(n178), .ZN(shiftedA_29__32_) );
  NOR2_X1 U1558 ( .A1(n167), .A2(n178), .ZN(shiftedA_29__31_) );
  NOR2_X1 U1559 ( .A1(n168), .A2(n178), .ZN(shiftedA_29__30_) );
  NOR2_X1 U1560 ( .A1(n136), .A2(n178), .ZN(shiftedA_29__29_) );
  NOR2_X1 U1561 ( .A1(n138), .A2(n179), .ZN(shiftedA_28__63_) );
  NOR2_X1 U1562 ( .A1(n139), .A2(n179), .ZN(shiftedA_28__58_) );
  NOR2_X1 U1563 ( .A1(n140), .A2(n179), .ZN(shiftedA_28__57_) );
  NOR2_X1 U1564 ( .A1(n141), .A2(n179), .ZN(shiftedA_28__56_) );
  NOR2_X1 U1565 ( .A1(n142), .A2(n179), .ZN(shiftedA_28__55_) );
  NOR2_X1 U1566 ( .A1(n143), .A2(n179), .ZN(shiftedA_28__54_) );
  NOR2_X1 U1567 ( .A1(n144), .A2(n179), .ZN(shiftedA_28__53_) );
  NOR2_X1 U1568 ( .A1(n145), .A2(n179), .ZN(shiftedA_28__52_) );
  NOR2_X1 U1569 ( .A1(n146), .A2(n179), .ZN(shiftedA_28__51_) );
  NOR2_X1 U1570 ( .A1(n147), .A2(n179), .ZN(shiftedA_28__50_) );
  NOR2_X1 U1571 ( .A1(n148), .A2(n179), .ZN(shiftedA_28__49_) );
  NOR2_X1 U1572 ( .A1(n149), .A2(n179), .ZN(shiftedA_28__48_) );
  NOR2_X1 U1573 ( .A1(n150), .A2(n179), .ZN(shiftedA_28__47_) );
  NOR2_X1 U1574 ( .A1(n151), .A2(n179), .ZN(shiftedA_28__46_) );
  NOR2_X1 U1575 ( .A1(n152), .A2(n179), .ZN(shiftedA_28__45_) );
  NOR2_X1 U1576 ( .A1(n153), .A2(n179), .ZN(shiftedA_28__44_) );
  NOR2_X1 U1577 ( .A1(n154), .A2(n179), .ZN(shiftedA_28__43_) );
  NOR2_X1 U1578 ( .A1(n155), .A2(n179), .ZN(shiftedA_28__42_) );
  NOR2_X1 U1579 ( .A1(n156), .A2(n179), .ZN(shiftedA_28__41_) );
  NOR2_X1 U1580 ( .A1(n157), .A2(n179), .ZN(shiftedA_28__40_) );
  NOR2_X1 U1581 ( .A1(n158), .A2(n179), .ZN(shiftedA_28__39_) );
  NOR2_X1 U1582 ( .A1(n159), .A2(n179), .ZN(shiftedA_28__38_) );
  NOR2_X1 U1583 ( .A1(n160), .A2(n179), .ZN(shiftedA_28__37_) );
  NOR2_X1 U1584 ( .A1(n161), .A2(n179), .ZN(shiftedA_28__36_) );
  NOR2_X1 U1585 ( .A1(n162), .A2(n179), .ZN(shiftedA_28__35_) );
  NOR2_X1 U1586 ( .A1(n163), .A2(n179), .ZN(shiftedA_28__34_) );
  NOR2_X1 U1587 ( .A1(n164), .A2(n179), .ZN(shiftedA_28__33_) );
  NOR2_X1 U1588 ( .A1(n165), .A2(n179), .ZN(shiftedA_28__32_) );
  NOR2_X1 U1589 ( .A1(n166), .A2(n179), .ZN(shiftedA_28__31_) );
  NOR2_X1 U1590 ( .A1(n167), .A2(n179), .ZN(shiftedA_28__30_) );
  NOR2_X1 U1591 ( .A1(n168), .A2(n179), .ZN(shiftedA_28__29_) );
  NOR2_X1 U1592 ( .A1(n136), .A2(n179), .ZN(shiftedA_28__28_) );
  NOR2_X1 U1593 ( .A1(n138), .A2(n180), .ZN(shiftedA_27__63_) );
  NOR2_X1 U1594 ( .A1(n139), .A2(n180), .ZN(shiftedA_27__57_) );
  NOR2_X1 U1595 ( .A1(n140), .A2(n180), .ZN(shiftedA_27__56_) );
  NOR2_X1 U1596 ( .A1(n141), .A2(n180), .ZN(shiftedA_27__55_) );
  NOR2_X1 U1597 ( .A1(n142), .A2(n180), .ZN(shiftedA_27__54_) );
  NOR2_X1 U1598 ( .A1(n143), .A2(n180), .ZN(shiftedA_27__53_) );
  NOR2_X1 U1599 ( .A1(n144), .A2(n180), .ZN(shiftedA_27__52_) );
  NOR2_X1 U1600 ( .A1(n145), .A2(n180), .ZN(shiftedA_27__51_) );
  NOR2_X1 U1601 ( .A1(n146), .A2(n180), .ZN(shiftedA_27__50_) );
  NOR2_X1 U1602 ( .A1(n147), .A2(n180), .ZN(shiftedA_27__49_) );
  NOR2_X1 U1603 ( .A1(n148), .A2(n180), .ZN(shiftedA_27__48_) );
  NOR2_X1 U1604 ( .A1(n149), .A2(n180), .ZN(shiftedA_27__47_) );
  NOR2_X1 U1605 ( .A1(n150), .A2(n180), .ZN(shiftedA_27__46_) );
  NOR2_X1 U1606 ( .A1(n151), .A2(n180), .ZN(shiftedA_27__45_) );
  NOR2_X1 U1607 ( .A1(n152), .A2(n180), .ZN(shiftedA_27__44_) );
  NOR2_X1 U1608 ( .A1(n153), .A2(n180), .ZN(shiftedA_27__43_) );
  NOR2_X1 U1609 ( .A1(n154), .A2(n180), .ZN(shiftedA_27__42_) );
  NOR2_X1 U1610 ( .A1(n155), .A2(n180), .ZN(shiftedA_27__41_) );
  NOR2_X1 U1611 ( .A1(n156), .A2(n180), .ZN(shiftedA_27__40_) );
  NOR2_X1 U1612 ( .A1(n157), .A2(n180), .ZN(shiftedA_27__39_) );
  NOR2_X1 U1613 ( .A1(n158), .A2(n180), .ZN(shiftedA_27__38_) );
  NOR2_X1 U1614 ( .A1(n159), .A2(n180), .ZN(shiftedA_27__37_) );
  NOR2_X1 U1615 ( .A1(n160), .A2(n180), .ZN(shiftedA_27__36_) );
  NOR2_X1 U1616 ( .A1(n161), .A2(n180), .ZN(shiftedA_27__35_) );
  NOR2_X1 U1617 ( .A1(n162), .A2(n180), .ZN(shiftedA_27__34_) );
  NOR2_X1 U1618 ( .A1(n163), .A2(n180), .ZN(shiftedA_27__33_) );
  NOR2_X1 U1619 ( .A1(n164), .A2(n180), .ZN(shiftedA_27__32_) );
  NOR2_X1 U1620 ( .A1(n165), .A2(n180), .ZN(shiftedA_27__31_) );
  NOR2_X1 U1621 ( .A1(n166), .A2(n180), .ZN(shiftedA_27__30_) );
  NOR2_X1 U1622 ( .A1(n167), .A2(n180), .ZN(shiftedA_27__29_) );
  NOR2_X1 U1623 ( .A1(n168), .A2(n180), .ZN(shiftedA_27__28_) );
  NOR2_X1 U1624 ( .A1(n136), .A2(n180), .ZN(shiftedA_27__27_) );
  NOR2_X1 U1625 ( .A1(n139), .A2(n181), .ZN(shiftedA_26__56_) );
  NOR2_X1 U1626 ( .A1(n140), .A2(n181), .ZN(shiftedA_26__55_) );
  NOR2_X1 U1627 ( .A1(n141), .A2(n181), .ZN(shiftedA_26__54_) );
  NOR2_X1 U1628 ( .A1(n142), .A2(n181), .ZN(shiftedA_26__53_) );
  NOR2_X1 U1629 ( .A1(n143), .A2(n181), .ZN(shiftedA_26__52_) );
  NOR2_X1 U1630 ( .A1(n144), .A2(n181), .ZN(shiftedA_26__51_) );
  NOR2_X1 U1631 ( .A1(n145), .A2(n181), .ZN(shiftedA_26__50_) );
  NOR2_X1 U1632 ( .A1(n146), .A2(n181), .ZN(shiftedA_26__49_) );
  NOR2_X1 U1633 ( .A1(n147), .A2(n181), .ZN(shiftedA_26__48_) );
  NOR2_X1 U1634 ( .A1(n148), .A2(n181), .ZN(shiftedA_26__47_) );
  NOR2_X1 U1635 ( .A1(n149), .A2(n181), .ZN(shiftedA_26__46_) );
  NOR2_X1 U1636 ( .A1(n150), .A2(n181), .ZN(shiftedA_26__45_) );
  NOR2_X1 U1637 ( .A1(n151), .A2(n181), .ZN(shiftedA_26__44_) );
  NOR2_X1 U1638 ( .A1(n152), .A2(n181), .ZN(shiftedA_26__43_) );
  NOR2_X1 U1639 ( .A1(n153), .A2(n181), .ZN(shiftedA_26__42_) );
  NOR2_X1 U1640 ( .A1(n154), .A2(n181), .ZN(shiftedA_26__41_) );
  NOR2_X1 U1641 ( .A1(n155), .A2(n181), .ZN(shiftedA_26__40_) );
  NOR2_X1 U1642 ( .A1(n156), .A2(n181), .ZN(shiftedA_26__39_) );
  NOR2_X1 U1643 ( .A1(n157), .A2(n181), .ZN(shiftedA_26__38_) );
  NOR2_X1 U1644 ( .A1(n158), .A2(n181), .ZN(shiftedA_26__37_) );
  NOR2_X1 U1645 ( .A1(n159), .A2(n181), .ZN(shiftedA_26__36_) );
  NOR2_X1 U1646 ( .A1(n160), .A2(n181), .ZN(shiftedA_26__35_) );
  NOR2_X1 U1647 ( .A1(n161), .A2(n181), .ZN(shiftedA_26__34_) );
  NOR2_X1 U1648 ( .A1(n162), .A2(n181), .ZN(shiftedA_26__33_) );
  NOR2_X1 U1649 ( .A1(n163), .A2(n181), .ZN(shiftedA_26__32_) );
  NOR2_X1 U1650 ( .A1(n164), .A2(n181), .ZN(shiftedA_26__31_) );
  NOR2_X1 U1651 ( .A1(n165), .A2(n181), .ZN(shiftedA_26__30_) );
  NOR2_X1 U1652 ( .A1(n166), .A2(n181), .ZN(shiftedA_26__29_) );
  NOR2_X1 U1653 ( .A1(n167), .A2(n181), .ZN(shiftedA_26__28_) );
  NOR2_X1 U1654 ( .A1(n168), .A2(n181), .ZN(shiftedA_26__27_) );
  NOR2_X1 U1655 ( .A1(n136), .A2(n181), .ZN(shiftedA_26__26_) );
  NOR2_X1 U1656 ( .A1(n139), .A2(n182), .ZN(shiftedA_25__55_) );
  NOR2_X1 U1657 ( .A1(n140), .A2(n182), .ZN(shiftedA_25__54_) );
  NOR2_X1 U1658 ( .A1(n141), .A2(n182), .ZN(shiftedA_25__53_) );
  NOR2_X1 U1659 ( .A1(n142), .A2(n182), .ZN(shiftedA_25__52_) );
  NOR2_X1 U1660 ( .A1(n143), .A2(n182), .ZN(shiftedA_25__51_) );
  NOR2_X1 U1661 ( .A1(n144), .A2(n182), .ZN(shiftedA_25__50_) );
  NOR2_X1 U1662 ( .A1(n145), .A2(n182), .ZN(shiftedA_25__49_) );
  NOR2_X1 U1663 ( .A1(n146), .A2(n182), .ZN(shiftedA_25__48_) );
  NOR2_X1 U1664 ( .A1(n147), .A2(n182), .ZN(shiftedA_25__47_) );
  NOR2_X1 U1665 ( .A1(n148), .A2(n182), .ZN(shiftedA_25__46_) );
  NOR2_X1 U1666 ( .A1(n149), .A2(n182), .ZN(shiftedA_25__45_) );
  NOR2_X1 U1667 ( .A1(n150), .A2(n182), .ZN(shiftedA_25__44_) );
  NOR2_X1 U1668 ( .A1(n151), .A2(n182), .ZN(shiftedA_25__43_) );
  NOR2_X1 U1669 ( .A1(n152), .A2(n182), .ZN(shiftedA_25__42_) );
  NOR2_X1 U1670 ( .A1(n153), .A2(n182), .ZN(shiftedA_25__41_) );
  NOR2_X1 U1671 ( .A1(n154), .A2(n182), .ZN(shiftedA_25__40_) );
  NOR2_X1 U1672 ( .A1(n155), .A2(n182), .ZN(shiftedA_25__39_) );
  NOR2_X1 U1673 ( .A1(n156), .A2(n182), .ZN(shiftedA_25__38_) );
  NOR2_X1 U1674 ( .A1(n157), .A2(n182), .ZN(shiftedA_25__37_) );
  NOR2_X1 U1675 ( .A1(n158), .A2(n182), .ZN(shiftedA_25__36_) );
  NOR2_X1 U1676 ( .A1(n159), .A2(n182), .ZN(shiftedA_25__35_) );
  NOR2_X1 U1677 ( .A1(n160), .A2(n182), .ZN(shiftedA_25__34_) );
  NOR2_X1 U1678 ( .A1(n161), .A2(n182), .ZN(shiftedA_25__33_) );
  NOR2_X1 U1679 ( .A1(n162), .A2(n182), .ZN(shiftedA_25__32_) );
  NOR2_X1 U1680 ( .A1(n163), .A2(n182), .ZN(shiftedA_25__31_) );
  NOR2_X1 U1681 ( .A1(n164), .A2(n182), .ZN(shiftedA_25__30_) );
  NOR2_X1 U1682 ( .A1(n165), .A2(n182), .ZN(shiftedA_25__29_) );
  NOR2_X1 U1683 ( .A1(n166), .A2(n182), .ZN(shiftedA_25__28_) );
  NOR2_X1 U1684 ( .A1(n167), .A2(n182), .ZN(shiftedA_25__27_) );
  NOR2_X1 U1685 ( .A1(n168), .A2(n182), .ZN(shiftedA_25__26_) );
  NOR2_X1 U1686 ( .A1(n136), .A2(n182), .ZN(shiftedA_25__25_) );
  NOR2_X1 U1687 ( .A1(n139), .A2(n183), .ZN(shiftedA_24__54_) );
  NOR2_X1 U1688 ( .A1(n140), .A2(n183), .ZN(shiftedA_24__53_) );
  NOR2_X1 U1689 ( .A1(n141), .A2(n183), .ZN(shiftedA_24__52_) );
  NOR2_X1 U1690 ( .A1(n142), .A2(n183), .ZN(shiftedA_24__51_) );
  NOR2_X1 U1691 ( .A1(n143), .A2(n183), .ZN(shiftedA_24__50_) );
  NOR2_X1 U1692 ( .A1(n144), .A2(n183), .ZN(shiftedA_24__49_) );
  NOR2_X1 U1693 ( .A1(n145), .A2(n183), .ZN(shiftedA_24__48_) );
  NOR2_X1 U1694 ( .A1(n146), .A2(n183), .ZN(shiftedA_24__47_) );
  NOR2_X1 U1695 ( .A1(n147), .A2(n183), .ZN(shiftedA_24__46_) );
  NOR2_X1 U1696 ( .A1(n148), .A2(n183), .ZN(shiftedA_24__45_) );
  NOR2_X1 U1697 ( .A1(n149), .A2(n183), .ZN(shiftedA_24__44_) );
  NOR2_X1 U1698 ( .A1(n150), .A2(n183), .ZN(shiftedA_24__43_) );
  NOR2_X1 U1699 ( .A1(n151), .A2(n183), .ZN(shiftedA_24__42_) );
  NOR2_X1 U1700 ( .A1(n152), .A2(n183), .ZN(shiftedA_24__41_) );
  NOR2_X1 U1701 ( .A1(n153), .A2(n183), .ZN(shiftedA_24__40_) );
  NOR2_X1 U1702 ( .A1(n154), .A2(n183), .ZN(shiftedA_24__39_) );
  NOR2_X1 U1703 ( .A1(n155), .A2(n183), .ZN(shiftedA_24__38_) );
  NOR2_X1 U1704 ( .A1(n156), .A2(n183), .ZN(shiftedA_24__37_) );
  NOR2_X1 U1705 ( .A1(n157), .A2(n183), .ZN(shiftedA_24__36_) );
  NOR2_X1 U1706 ( .A1(n158), .A2(n183), .ZN(shiftedA_24__35_) );
  NOR2_X1 U1707 ( .A1(n159), .A2(n183), .ZN(shiftedA_24__34_) );
  NOR2_X1 U1708 ( .A1(n160), .A2(n183), .ZN(shiftedA_24__33_) );
  NOR2_X1 U1709 ( .A1(n161), .A2(n183), .ZN(shiftedA_24__32_) );
  NOR2_X1 U1710 ( .A1(n162), .A2(n183), .ZN(shiftedA_24__31_) );
  NOR2_X1 U1711 ( .A1(n163), .A2(n183), .ZN(shiftedA_24__30_) );
  NOR2_X1 U1712 ( .A1(n164), .A2(n183), .ZN(shiftedA_24__29_) );
  NOR2_X1 U1713 ( .A1(n165), .A2(n183), .ZN(shiftedA_24__28_) );
  NOR2_X1 U1714 ( .A1(n166), .A2(n183), .ZN(shiftedA_24__27_) );
  NOR2_X1 U1715 ( .A1(n167), .A2(n183), .ZN(shiftedA_24__26_) );
  NOR2_X1 U1716 ( .A1(n168), .A2(n183), .ZN(shiftedA_24__25_) );
  NOR2_X1 U1717 ( .A1(n136), .A2(n183), .ZN(shiftedA_24__24_) );
  NOR2_X1 U1718 ( .A1(n139), .A2(n184), .ZN(shiftedA_23__53_) );
  NOR2_X1 U1719 ( .A1(n140), .A2(n184), .ZN(shiftedA_23__52_) );
  NOR2_X1 U1720 ( .A1(n141), .A2(n184), .ZN(shiftedA_23__51_) );
  NOR2_X1 U1721 ( .A1(n142), .A2(n184), .ZN(shiftedA_23__50_) );
  NOR2_X1 U1722 ( .A1(n143), .A2(n184), .ZN(shiftedA_23__49_) );
  NOR2_X1 U1723 ( .A1(n144), .A2(n184), .ZN(shiftedA_23__48_) );
  NOR2_X1 U1724 ( .A1(n145), .A2(n184), .ZN(shiftedA_23__47_) );
  NOR2_X1 U1725 ( .A1(n146), .A2(n184), .ZN(shiftedA_23__46_) );
  NOR2_X1 U1726 ( .A1(n147), .A2(n184), .ZN(shiftedA_23__45_) );
  NOR2_X1 U1727 ( .A1(n148), .A2(n184), .ZN(shiftedA_23__44_) );
  NOR2_X1 U1728 ( .A1(n149), .A2(n184), .ZN(shiftedA_23__43_) );
  NOR2_X1 U1729 ( .A1(n150), .A2(n184), .ZN(shiftedA_23__42_) );
  NOR2_X1 U1730 ( .A1(n151), .A2(n184), .ZN(shiftedA_23__41_) );
  NOR2_X1 U1731 ( .A1(n152), .A2(n184), .ZN(shiftedA_23__40_) );
  NOR2_X1 U1732 ( .A1(n153), .A2(n184), .ZN(shiftedA_23__39_) );
  NOR2_X1 U1733 ( .A1(n154), .A2(n184), .ZN(shiftedA_23__38_) );
  NOR2_X1 U1734 ( .A1(n155), .A2(n184), .ZN(shiftedA_23__37_) );
  NOR2_X1 U1735 ( .A1(n156), .A2(n184), .ZN(shiftedA_23__36_) );
  NOR2_X1 U1736 ( .A1(n157), .A2(n184), .ZN(shiftedA_23__35_) );
  NOR2_X1 U1737 ( .A1(n158), .A2(n184), .ZN(shiftedA_23__34_) );
  NOR2_X1 U1738 ( .A1(n159), .A2(n184), .ZN(shiftedA_23__33_) );
  NOR2_X1 U1739 ( .A1(n160), .A2(n184), .ZN(shiftedA_23__32_) );
  NOR2_X1 U1740 ( .A1(n161), .A2(n184), .ZN(shiftedA_23__31_) );
  NOR2_X1 U1741 ( .A1(n162), .A2(n184), .ZN(shiftedA_23__30_) );
  NOR2_X1 U1742 ( .A1(n163), .A2(n184), .ZN(shiftedA_23__29_) );
  NOR2_X1 U1743 ( .A1(n164), .A2(n184), .ZN(shiftedA_23__28_) );
  NOR2_X1 U1744 ( .A1(n165), .A2(n184), .ZN(shiftedA_23__27_) );
  NOR2_X1 U1745 ( .A1(n166), .A2(n184), .ZN(shiftedA_23__26_) );
  NOR2_X1 U1746 ( .A1(n167), .A2(n184), .ZN(shiftedA_23__25_) );
  NOR2_X1 U1747 ( .A1(n168), .A2(n184), .ZN(shiftedA_23__24_) );
  NOR2_X1 U1748 ( .A1(n136), .A2(n184), .ZN(shiftedA_23__23_) );
  NOR2_X1 U1749 ( .A1(n139), .A2(n185), .ZN(shiftedA_22__52_) );
  NOR2_X1 U1750 ( .A1(n140), .A2(n185), .ZN(shiftedA_22__51_) );
  NOR2_X1 U1751 ( .A1(n141), .A2(n185), .ZN(shiftedA_22__50_) );
  NOR2_X1 U1752 ( .A1(n142), .A2(n185), .ZN(shiftedA_22__49_) );
  NOR2_X1 U1753 ( .A1(n143), .A2(n185), .ZN(shiftedA_22__48_) );
  NOR2_X1 U1754 ( .A1(n144), .A2(n185), .ZN(shiftedA_22__47_) );
  NOR2_X1 U1755 ( .A1(n145), .A2(n185), .ZN(shiftedA_22__46_) );
  NOR2_X1 U1756 ( .A1(n146), .A2(n185), .ZN(shiftedA_22__45_) );
  NOR2_X1 U1757 ( .A1(n147), .A2(n185), .ZN(shiftedA_22__44_) );
  NOR2_X1 U1758 ( .A1(n148), .A2(n185), .ZN(shiftedA_22__43_) );
  NOR2_X1 U1759 ( .A1(n149), .A2(n185), .ZN(shiftedA_22__42_) );
  NOR2_X1 U1760 ( .A1(n150), .A2(n185), .ZN(shiftedA_22__41_) );
  NOR2_X1 U1761 ( .A1(n151), .A2(n185), .ZN(shiftedA_22__40_) );
  NOR2_X1 U1762 ( .A1(n152), .A2(n185), .ZN(shiftedA_22__39_) );
  NOR2_X1 U1763 ( .A1(n153), .A2(n185), .ZN(shiftedA_22__38_) );
  NOR2_X1 U1764 ( .A1(n154), .A2(n185), .ZN(shiftedA_22__37_) );
  NOR2_X1 U1765 ( .A1(n155), .A2(n185), .ZN(shiftedA_22__36_) );
  NOR2_X1 U1766 ( .A1(n156), .A2(n185), .ZN(shiftedA_22__35_) );
  NOR2_X1 U1767 ( .A1(n157), .A2(n185), .ZN(shiftedA_22__34_) );
  NOR2_X1 U1768 ( .A1(n158), .A2(n185), .ZN(shiftedA_22__33_) );
  NOR2_X1 U1769 ( .A1(n159), .A2(n185), .ZN(shiftedA_22__32_) );
  NOR2_X1 U1770 ( .A1(n160), .A2(n185), .ZN(shiftedA_22__31_) );
  NOR2_X1 U1771 ( .A1(n161), .A2(n185), .ZN(shiftedA_22__30_) );
  NOR2_X1 U1772 ( .A1(n162), .A2(n185), .ZN(shiftedA_22__29_) );
  NOR2_X1 U1773 ( .A1(n163), .A2(n185), .ZN(shiftedA_22__28_) );
  NOR2_X1 U1774 ( .A1(n164), .A2(n185), .ZN(shiftedA_22__27_) );
  NOR2_X1 U1775 ( .A1(n165), .A2(n185), .ZN(shiftedA_22__26_) );
  NOR2_X1 U1776 ( .A1(n166), .A2(n185), .ZN(shiftedA_22__25_) );
  NOR2_X1 U1777 ( .A1(n167), .A2(n185), .ZN(shiftedA_22__24_) );
  NOR2_X1 U1778 ( .A1(n168), .A2(n185), .ZN(shiftedA_22__23_) );
  NOR2_X1 U1779 ( .A1(n136), .A2(n185), .ZN(shiftedA_22__22_) );
  NOR2_X1 U1780 ( .A1(n139), .A2(n186), .ZN(shiftedA_21__51_) );
  NOR2_X1 U1781 ( .A1(n140), .A2(n186), .ZN(shiftedA_21__50_) );
  NOR2_X1 U1782 ( .A1(n141), .A2(n186), .ZN(shiftedA_21__49_) );
  NOR2_X1 U1783 ( .A1(n142), .A2(n186), .ZN(shiftedA_21__48_) );
  NOR2_X1 U1784 ( .A1(n143), .A2(n186), .ZN(shiftedA_21__47_) );
  NOR2_X1 U1785 ( .A1(n144), .A2(n186), .ZN(shiftedA_21__46_) );
  NOR2_X1 U1786 ( .A1(n145), .A2(n186), .ZN(shiftedA_21__45_) );
  NOR2_X1 U1787 ( .A1(n146), .A2(n186), .ZN(shiftedA_21__44_) );
  NOR2_X1 U1788 ( .A1(n147), .A2(n186), .ZN(shiftedA_21__43_) );
  NOR2_X1 U1789 ( .A1(n148), .A2(n186), .ZN(shiftedA_21__42_) );
  NOR2_X1 U1790 ( .A1(n149), .A2(n186), .ZN(shiftedA_21__41_) );
  NOR2_X1 U1791 ( .A1(n150), .A2(n186), .ZN(shiftedA_21__40_) );
  NOR2_X1 U1792 ( .A1(n151), .A2(n186), .ZN(shiftedA_21__39_) );
  NOR2_X1 U1793 ( .A1(n152), .A2(n186), .ZN(shiftedA_21__38_) );
  NOR2_X1 U1794 ( .A1(n153), .A2(n186), .ZN(shiftedA_21__37_) );
  NOR2_X1 U1795 ( .A1(n154), .A2(n186), .ZN(shiftedA_21__36_) );
  NOR2_X1 U1796 ( .A1(n155), .A2(n186), .ZN(shiftedA_21__35_) );
  NOR2_X1 U1797 ( .A1(n156), .A2(n186), .ZN(shiftedA_21__34_) );
  NOR2_X1 U1798 ( .A1(n157), .A2(n186), .ZN(shiftedA_21__33_) );
  NOR2_X1 U1799 ( .A1(n158), .A2(n186), .ZN(shiftedA_21__32_) );
  NOR2_X1 U1800 ( .A1(n159), .A2(n186), .ZN(shiftedA_21__31_) );
  NOR2_X1 U1801 ( .A1(n160), .A2(n186), .ZN(shiftedA_21__30_) );
  NOR2_X1 U1802 ( .A1(n161), .A2(n186), .ZN(shiftedA_21__29_) );
  NOR2_X1 U1803 ( .A1(n162), .A2(n186), .ZN(shiftedA_21__28_) );
  NOR2_X1 U1804 ( .A1(n163), .A2(n186), .ZN(shiftedA_21__27_) );
  NOR2_X1 U1805 ( .A1(n164), .A2(n186), .ZN(shiftedA_21__26_) );
  NOR2_X1 U1806 ( .A1(n165), .A2(n186), .ZN(shiftedA_21__25_) );
  NOR2_X1 U1807 ( .A1(n166), .A2(n186), .ZN(shiftedA_21__24_) );
  NOR2_X1 U1808 ( .A1(n167), .A2(n186), .ZN(shiftedA_21__23_) );
  NOR2_X1 U1809 ( .A1(n168), .A2(n186), .ZN(shiftedA_21__22_) );
  NOR2_X1 U1810 ( .A1(n136), .A2(n186), .ZN(shiftedA_21__21_) );
  NOR2_X1 U1811 ( .A1(n139), .A2(n187), .ZN(shiftedA_20__50_) );
  NOR2_X1 U1812 ( .A1(n140), .A2(n187), .ZN(shiftedA_20__49_) );
  NOR2_X1 U1813 ( .A1(n141), .A2(n187), .ZN(shiftedA_20__48_) );
  NOR2_X1 U1814 ( .A1(n142), .A2(n187), .ZN(shiftedA_20__47_) );
  NOR2_X1 U1815 ( .A1(n143), .A2(n187), .ZN(shiftedA_20__46_) );
  NOR2_X1 U1816 ( .A1(n144), .A2(n187), .ZN(shiftedA_20__45_) );
  NOR2_X1 U1817 ( .A1(n145), .A2(n187), .ZN(shiftedA_20__44_) );
  NOR2_X1 U1818 ( .A1(n146), .A2(n187), .ZN(shiftedA_20__43_) );
  NOR2_X1 U1819 ( .A1(n147), .A2(n187), .ZN(shiftedA_20__42_) );
  NOR2_X1 U1820 ( .A1(n148), .A2(n187), .ZN(shiftedA_20__41_) );
  NOR2_X1 U1821 ( .A1(n149), .A2(n187), .ZN(shiftedA_20__40_) );
  NOR2_X1 U1822 ( .A1(n150), .A2(n187), .ZN(shiftedA_20__39_) );
  NOR2_X1 U1823 ( .A1(n151), .A2(n187), .ZN(shiftedA_20__38_) );
  NOR2_X1 U1824 ( .A1(n152), .A2(n187), .ZN(shiftedA_20__37_) );
  NOR2_X1 U1825 ( .A1(n153), .A2(n187), .ZN(shiftedA_20__36_) );
  NOR2_X1 U1826 ( .A1(n154), .A2(n187), .ZN(shiftedA_20__35_) );
  NOR2_X1 U1827 ( .A1(n155), .A2(n187), .ZN(shiftedA_20__34_) );
  NOR2_X1 U1828 ( .A1(n156), .A2(n187), .ZN(shiftedA_20__33_) );
  NOR2_X1 U1829 ( .A1(n157), .A2(n187), .ZN(shiftedA_20__32_) );
  NOR2_X1 U1830 ( .A1(n158), .A2(n187), .ZN(shiftedA_20__31_) );
  NOR2_X1 U1831 ( .A1(n159), .A2(n187), .ZN(shiftedA_20__30_) );
  NOR2_X1 U1832 ( .A1(n160), .A2(n187), .ZN(shiftedA_20__29_) );
  NOR2_X1 U1833 ( .A1(n161), .A2(n187), .ZN(shiftedA_20__28_) );
  NOR2_X1 U1834 ( .A1(n162), .A2(n187), .ZN(shiftedA_20__27_) );
  NOR2_X1 U1835 ( .A1(n163), .A2(n187), .ZN(shiftedA_20__26_) );
  NOR2_X1 U1836 ( .A1(n164), .A2(n187), .ZN(shiftedA_20__25_) );
  NOR2_X1 U1837 ( .A1(n165), .A2(n187), .ZN(shiftedA_20__24_) );
  NOR2_X1 U1838 ( .A1(n166), .A2(n187), .ZN(shiftedA_20__23_) );
  NOR2_X1 U1839 ( .A1(n167), .A2(n187), .ZN(shiftedA_20__22_) );
  NOR2_X1 U1840 ( .A1(n168), .A2(n187), .ZN(shiftedA_20__21_) );
  NOR2_X1 U1841 ( .A1(n136), .A2(n187), .ZN(shiftedA_20__20_) );
  NOR2_X1 U1842 ( .A1(n161), .A2(n188), .ZN(shiftedA_1__9_) );
  NOR2_X1 U1843 ( .A1(n162), .A2(n188), .ZN(shiftedA_1__8_) );
  NOR2_X1 U1844 ( .A1(n163), .A2(n188), .ZN(shiftedA_1__7_) );
  NOR2_X1 U1845 ( .A1(n164), .A2(n188), .ZN(shiftedA_1__6_) );
  NOR2_X1 U1846 ( .A1(n165), .A2(n188), .ZN(shiftedA_1__5_) );
  NOR2_X1 U1847 ( .A1(n166), .A2(n188), .ZN(shiftedA_1__4_) );
  NOR2_X1 U1848 ( .A1(n167), .A2(n188), .ZN(shiftedA_1__3_) );
  NOR2_X1 U1849 ( .A1(n139), .A2(n188), .ZN(shiftedA_1__31_) );
  NOR2_X1 U1850 ( .A1(n140), .A2(n188), .ZN(shiftedA_1__30_) );
  NOR2_X1 U1851 ( .A1(n168), .A2(n188), .ZN(shiftedA_1__2_) );
  NOR2_X1 U1852 ( .A1(n141), .A2(n188), .ZN(shiftedA_1__29_) );
  NOR2_X1 U1853 ( .A1(n142), .A2(n188), .ZN(shiftedA_1__28_) );
  NOR2_X1 U1854 ( .A1(n143), .A2(n188), .ZN(shiftedA_1__27_) );
  NOR2_X1 U1855 ( .A1(n144), .A2(n188), .ZN(shiftedA_1__26_) );
  NOR2_X1 U1856 ( .A1(n145), .A2(n188), .ZN(shiftedA_1__25_) );
  NOR2_X1 U1857 ( .A1(n146), .A2(n188), .ZN(shiftedA_1__24_) );
  NOR2_X1 U1858 ( .A1(n147), .A2(n188), .ZN(shiftedA_1__23_) );
  NOR2_X1 U1859 ( .A1(n148), .A2(n188), .ZN(shiftedA_1__22_) );
  NOR2_X1 U1860 ( .A1(n149), .A2(n188), .ZN(shiftedA_1__21_) );
  NOR2_X1 U1861 ( .A1(n150), .A2(n188), .ZN(shiftedA_1__20_) );
  NOR2_X1 U1862 ( .A1(n136), .A2(n188), .ZN(shiftedA_1__1_) );
  NOR2_X1 U1863 ( .A1(n151), .A2(n188), .ZN(shiftedA_1__19_) );
  NOR2_X1 U1864 ( .A1(n152), .A2(n188), .ZN(shiftedA_1__18_) );
  NOR2_X1 U1865 ( .A1(n153), .A2(n188), .ZN(shiftedA_1__17_) );
  NOR2_X1 U1866 ( .A1(n154), .A2(n188), .ZN(shiftedA_1__16_) );
  NOR2_X1 U1867 ( .A1(n155), .A2(n188), .ZN(shiftedA_1__15_) );
  NOR2_X1 U1868 ( .A1(n156), .A2(n188), .ZN(shiftedA_1__14_) );
  NOR2_X1 U1869 ( .A1(n157), .A2(n188), .ZN(shiftedA_1__13_) );
  NOR2_X1 U1870 ( .A1(n158), .A2(n188), .ZN(shiftedA_1__12_) );
  NOR2_X1 U1871 ( .A1(n159), .A2(n188), .ZN(shiftedA_1__11_) );
  NOR2_X1 U1872 ( .A1(n160), .A2(n188), .ZN(shiftedA_1__10_) );
  NOR2_X1 U1873 ( .A1(n139), .A2(n189), .ZN(shiftedA_19__49_) );
  NOR2_X1 U1874 ( .A1(n140), .A2(n189), .ZN(shiftedA_19__48_) );
  NOR2_X1 U1875 ( .A1(n141), .A2(n189), .ZN(shiftedA_19__47_) );
  NOR2_X1 U1876 ( .A1(n142), .A2(n189), .ZN(shiftedA_19__46_) );
  NOR2_X1 U1877 ( .A1(n143), .A2(n189), .ZN(shiftedA_19__45_) );
  NOR2_X1 U1878 ( .A1(n144), .A2(n189), .ZN(shiftedA_19__44_) );
  NOR2_X1 U1879 ( .A1(n145), .A2(n189), .ZN(shiftedA_19__43_) );
  NOR2_X1 U1880 ( .A1(n146), .A2(n189), .ZN(shiftedA_19__42_) );
  NOR2_X1 U1881 ( .A1(n147), .A2(n189), .ZN(shiftedA_19__41_) );
  NOR2_X1 U1882 ( .A1(n148), .A2(n189), .ZN(shiftedA_19__40_) );
  NOR2_X1 U1883 ( .A1(n149), .A2(n189), .ZN(shiftedA_19__39_) );
  NOR2_X1 U1884 ( .A1(n150), .A2(n189), .ZN(shiftedA_19__38_) );
  NOR2_X1 U1885 ( .A1(n151), .A2(n189), .ZN(shiftedA_19__37_) );
  NOR2_X1 U1886 ( .A1(n152), .A2(n189), .ZN(shiftedA_19__36_) );
  NOR2_X1 U1887 ( .A1(n153), .A2(n189), .ZN(shiftedA_19__35_) );
  NOR2_X1 U1888 ( .A1(n154), .A2(n189), .ZN(shiftedA_19__34_) );
  NOR2_X1 U1889 ( .A1(n155), .A2(n189), .ZN(shiftedA_19__33_) );
  NOR2_X1 U1890 ( .A1(n156), .A2(n189), .ZN(shiftedA_19__32_) );
  NOR2_X1 U1891 ( .A1(n157), .A2(n189), .ZN(shiftedA_19__31_) );
  NOR2_X1 U1892 ( .A1(n158), .A2(n189), .ZN(shiftedA_19__30_) );
  NOR2_X1 U1893 ( .A1(n159), .A2(n189), .ZN(shiftedA_19__29_) );
  NOR2_X1 U1894 ( .A1(n160), .A2(n189), .ZN(shiftedA_19__28_) );
  NOR2_X1 U1895 ( .A1(n161), .A2(n189), .ZN(shiftedA_19__27_) );
  NOR2_X1 U1896 ( .A1(n162), .A2(n189), .ZN(shiftedA_19__26_) );
  NOR2_X1 U1897 ( .A1(n163), .A2(n189), .ZN(shiftedA_19__25_) );
  NOR2_X1 U1898 ( .A1(n164), .A2(n189), .ZN(shiftedA_19__24_) );
  NOR2_X1 U1899 ( .A1(n165), .A2(n189), .ZN(shiftedA_19__23_) );
  NOR2_X1 U1900 ( .A1(n166), .A2(n189), .ZN(shiftedA_19__22_) );
  NOR2_X1 U1901 ( .A1(n167), .A2(n189), .ZN(shiftedA_19__21_) );
  NOR2_X1 U1902 ( .A1(n168), .A2(n189), .ZN(shiftedA_19__20_) );
  NOR2_X1 U1903 ( .A1(n136), .A2(n189), .ZN(shiftedA_19__19_) );
  NOR2_X1 U1904 ( .A1(n139), .A2(n190), .ZN(shiftedA_18__48_) );
  NOR2_X1 U1905 ( .A1(n140), .A2(n190), .ZN(shiftedA_18__47_) );
  NOR2_X1 U1906 ( .A1(n141), .A2(n190), .ZN(shiftedA_18__46_) );
  NOR2_X1 U1907 ( .A1(n142), .A2(n190), .ZN(shiftedA_18__45_) );
  NOR2_X1 U1908 ( .A1(n143), .A2(n190), .ZN(shiftedA_18__44_) );
  NOR2_X1 U1909 ( .A1(n144), .A2(n190), .ZN(shiftedA_18__43_) );
  NOR2_X1 U1910 ( .A1(n145), .A2(n190), .ZN(shiftedA_18__42_) );
  NOR2_X1 U1911 ( .A1(n146), .A2(n190), .ZN(shiftedA_18__41_) );
  NOR2_X1 U1912 ( .A1(n147), .A2(n190), .ZN(shiftedA_18__40_) );
  NOR2_X1 U1913 ( .A1(n148), .A2(n190), .ZN(shiftedA_18__39_) );
  NOR2_X1 U1914 ( .A1(n149), .A2(n190), .ZN(shiftedA_18__38_) );
  NOR2_X1 U1915 ( .A1(n150), .A2(n190), .ZN(shiftedA_18__37_) );
  NOR2_X1 U1916 ( .A1(n151), .A2(n190), .ZN(shiftedA_18__36_) );
  NOR2_X1 U1917 ( .A1(n152), .A2(n190), .ZN(shiftedA_18__35_) );
  NOR2_X1 U1918 ( .A1(n153), .A2(n190), .ZN(shiftedA_18__34_) );
  NOR2_X1 U1919 ( .A1(n154), .A2(n190), .ZN(shiftedA_18__33_) );
  NOR2_X1 U1920 ( .A1(n155), .A2(n190), .ZN(shiftedA_18__32_) );
  NOR2_X1 U1921 ( .A1(n156), .A2(n190), .ZN(shiftedA_18__31_) );
  NOR2_X1 U1922 ( .A1(n157), .A2(n190), .ZN(shiftedA_18__30_) );
  NOR2_X1 U1923 ( .A1(n158), .A2(n190), .ZN(shiftedA_18__29_) );
  NOR2_X1 U1924 ( .A1(n159), .A2(n190), .ZN(shiftedA_18__28_) );
  NOR2_X1 U1925 ( .A1(n160), .A2(n190), .ZN(shiftedA_18__27_) );
  NOR2_X1 U1926 ( .A1(n161), .A2(n190), .ZN(shiftedA_18__26_) );
  NOR2_X1 U1927 ( .A1(n162), .A2(n190), .ZN(shiftedA_18__25_) );
  NOR2_X1 U1928 ( .A1(n163), .A2(n190), .ZN(shiftedA_18__24_) );
  NOR2_X1 U1929 ( .A1(n164), .A2(n190), .ZN(shiftedA_18__23_) );
  NOR2_X1 U1930 ( .A1(n165), .A2(n190), .ZN(shiftedA_18__22_) );
  NOR2_X1 U1931 ( .A1(n166), .A2(n190), .ZN(shiftedA_18__21_) );
  NOR2_X1 U1932 ( .A1(n167), .A2(n190), .ZN(shiftedA_18__20_) );
  NOR2_X1 U1933 ( .A1(n168), .A2(n190), .ZN(shiftedA_18__19_) );
  NOR2_X1 U1934 ( .A1(n136), .A2(n190), .ZN(shiftedA_18__18_) );
  NOR2_X1 U1935 ( .A1(n139), .A2(n191), .ZN(shiftedA_17__47_) );
  NOR2_X1 U1936 ( .A1(n140), .A2(n191), .ZN(shiftedA_17__46_) );
  NOR2_X1 U1937 ( .A1(n141), .A2(n191), .ZN(shiftedA_17__45_) );
  NOR2_X1 U1938 ( .A1(n142), .A2(n191), .ZN(shiftedA_17__44_) );
  NOR2_X1 U1939 ( .A1(n143), .A2(n191), .ZN(shiftedA_17__43_) );
  NOR2_X1 U1940 ( .A1(n144), .A2(n191), .ZN(shiftedA_17__42_) );
  NOR2_X1 U1941 ( .A1(n145), .A2(n191), .ZN(shiftedA_17__41_) );
  NOR2_X1 U1942 ( .A1(n146), .A2(n191), .ZN(shiftedA_17__40_) );
  NOR2_X1 U1943 ( .A1(n147), .A2(n191), .ZN(shiftedA_17__39_) );
  NOR2_X1 U1944 ( .A1(n148), .A2(n191), .ZN(shiftedA_17__38_) );
  NOR2_X1 U1945 ( .A1(n149), .A2(n191), .ZN(shiftedA_17__37_) );
  NOR2_X1 U1946 ( .A1(n150), .A2(n191), .ZN(shiftedA_17__36_) );
  NOR2_X1 U1947 ( .A1(n151), .A2(n191), .ZN(shiftedA_17__35_) );
  NOR2_X1 U1948 ( .A1(n152), .A2(n191), .ZN(shiftedA_17__34_) );
  NOR2_X1 U1949 ( .A1(n153), .A2(n191), .ZN(shiftedA_17__33_) );
  NOR2_X1 U1950 ( .A1(n154), .A2(n191), .ZN(shiftedA_17__32_) );
  NOR2_X1 U1951 ( .A1(n155), .A2(n191), .ZN(shiftedA_17__31_) );
  NOR2_X1 U1952 ( .A1(n156), .A2(n191), .ZN(shiftedA_17__30_) );
  NOR2_X1 U1953 ( .A1(n157), .A2(n191), .ZN(shiftedA_17__29_) );
  NOR2_X1 U1954 ( .A1(n158), .A2(n191), .ZN(shiftedA_17__28_) );
  NOR2_X1 U1955 ( .A1(n159), .A2(n191), .ZN(shiftedA_17__27_) );
  NOR2_X1 U1956 ( .A1(n160), .A2(n191), .ZN(shiftedA_17__26_) );
  NOR2_X1 U1957 ( .A1(n161), .A2(n191), .ZN(shiftedA_17__25_) );
  NOR2_X1 U1958 ( .A1(n162), .A2(n191), .ZN(shiftedA_17__24_) );
  NOR2_X1 U1959 ( .A1(n163), .A2(n191), .ZN(shiftedA_17__23_) );
  NOR2_X1 U1960 ( .A1(n164), .A2(n191), .ZN(shiftedA_17__22_) );
  NOR2_X1 U1961 ( .A1(n165), .A2(n191), .ZN(shiftedA_17__21_) );
  NOR2_X1 U1962 ( .A1(n166), .A2(n191), .ZN(shiftedA_17__20_) );
  NOR2_X1 U1963 ( .A1(n167), .A2(n191), .ZN(shiftedA_17__19_) );
  NOR2_X1 U1964 ( .A1(n168), .A2(n191), .ZN(shiftedA_17__18_) );
  NOR2_X1 U1965 ( .A1(n136), .A2(n191), .ZN(shiftedA_17__17_) );
  NOR2_X1 U1966 ( .A1(n139), .A2(n192), .ZN(shiftedA_16__46_) );
  NOR2_X1 U1967 ( .A1(n140), .A2(n192), .ZN(shiftedA_16__45_) );
  NOR2_X1 U1968 ( .A1(n141), .A2(n192), .ZN(shiftedA_16__44_) );
  NOR2_X1 U1969 ( .A1(n142), .A2(n192), .ZN(shiftedA_16__43_) );
  NOR2_X1 U1970 ( .A1(n143), .A2(n192), .ZN(shiftedA_16__42_) );
  NOR2_X1 U1971 ( .A1(n144), .A2(n192), .ZN(shiftedA_16__41_) );
  NOR2_X1 U1972 ( .A1(n145), .A2(n192), .ZN(shiftedA_16__40_) );
  NOR2_X1 U1973 ( .A1(n146), .A2(n192), .ZN(shiftedA_16__39_) );
  NOR2_X1 U1974 ( .A1(n147), .A2(n192), .ZN(shiftedA_16__38_) );
  NOR2_X1 U1975 ( .A1(n148), .A2(n192), .ZN(shiftedA_16__37_) );
  NOR2_X1 U1976 ( .A1(n149), .A2(n192), .ZN(shiftedA_16__36_) );
  NOR2_X1 U1977 ( .A1(n150), .A2(n192), .ZN(shiftedA_16__35_) );
  NOR2_X1 U1978 ( .A1(n151), .A2(n192), .ZN(shiftedA_16__34_) );
  NOR2_X1 U1979 ( .A1(n152), .A2(n192), .ZN(shiftedA_16__33_) );
  NOR2_X1 U1980 ( .A1(n153), .A2(n192), .ZN(shiftedA_16__32_) );
  NOR2_X1 U1981 ( .A1(n154), .A2(n192), .ZN(shiftedA_16__31_) );
  NOR2_X1 U1982 ( .A1(n155), .A2(n192), .ZN(shiftedA_16__30_) );
  NOR2_X1 U1983 ( .A1(n156), .A2(n192), .ZN(shiftedA_16__29_) );
  NOR2_X1 U1984 ( .A1(n157), .A2(n192), .ZN(shiftedA_16__28_) );
  NOR2_X1 U1985 ( .A1(n158), .A2(n192), .ZN(shiftedA_16__27_) );
  NOR2_X1 U1986 ( .A1(n159), .A2(n192), .ZN(shiftedA_16__26_) );
  NOR2_X1 U1987 ( .A1(n160), .A2(n192), .ZN(shiftedA_16__25_) );
  NOR2_X1 U1988 ( .A1(n161), .A2(n192), .ZN(shiftedA_16__24_) );
  NOR2_X1 U1989 ( .A1(n162), .A2(n192), .ZN(shiftedA_16__23_) );
  NOR2_X1 U1990 ( .A1(n163), .A2(n192), .ZN(shiftedA_16__22_) );
  NOR2_X1 U1991 ( .A1(n164), .A2(n192), .ZN(shiftedA_16__21_) );
  NOR2_X1 U1992 ( .A1(n165), .A2(n192), .ZN(shiftedA_16__20_) );
  NOR2_X1 U1993 ( .A1(n166), .A2(n192), .ZN(shiftedA_16__19_) );
  NOR2_X1 U1994 ( .A1(n167), .A2(n192), .ZN(shiftedA_16__18_) );
  NOR2_X1 U1995 ( .A1(n168), .A2(n192), .ZN(shiftedA_16__17_) );
  NOR2_X1 U1996 ( .A1(n136), .A2(n192), .ZN(shiftedA_16__16_) );
  NOR2_X1 U1997 ( .A1(n139), .A2(n193), .ZN(shiftedA_15__45_) );
  NOR2_X1 U1998 ( .A1(n140), .A2(n193), .ZN(shiftedA_15__44_) );
  NOR2_X1 U1999 ( .A1(n141), .A2(n193), .ZN(shiftedA_15__43_) );
  NOR2_X1 U2000 ( .A1(n142), .A2(n193), .ZN(shiftedA_15__42_) );
  NOR2_X1 U2001 ( .A1(n143), .A2(n193), .ZN(shiftedA_15__41_) );
  NOR2_X1 U2002 ( .A1(n144), .A2(n193), .ZN(shiftedA_15__40_) );
  NOR2_X1 U2003 ( .A1(n145), .A2(n193), .ZN(shiftedA_15__39_) );
  NOR2_X1 U2004 ( .A1(n146), .A2(n193), .ZN(shiftedA_15__38_) );
  NOR2_X1 U2005 ( .A1(n147), .A2(n193), .ZN(shiftedA_15__37_) );
  NOR2_X1 U2006 ( .A1(n148), .A2(n193), .ZN(shiftedA_15__36_) );
  NOR2_X1 U2007 ( .A1(n149), .A2(n193), .ZN(shiftedA_15__35_) );
  NOR2_X1 U2008 ( .A1(n150), .A2(n193), .ZN(shiftedA_15__34_) );
  NOR2_X1 U2009 ( .A1(n151), .A2(n193), .ZN(shiftedA_15__33_) );
  NOR2_X1 U2010 ( .A1(n152), .A2(n193), .ZN(shiftedA_15__32_) );
  NOR2_X1 U2011 ( .A1(n153), .A2(n193), .ZN(shiftedA_15__31_) );
  NOR2_X1 U2012 ( .A1(n154), .A2(n193), .ZN(shiftedA_15__30_) );
  NOR2_X1 U2013 ( .A1(n155), .A2(n193), .ZN(shiftedA_15__29_) );
  NOR2_X1 U2014 ( .A1(n156), .A2(n193), .ZN(shiftedA_15__28_) );
  NOR2_X1 U2015 ( .A1(n157), .A2(n193), .ZN(shiftedA_15__27_) );
  NOR2_X1 U2016 ( .A1(n158), .A2(n193), .ZN(shiftedA_15__26_) );
  NOR2_X1 U2017 ( .A1(n159), .A2(n193), .ZN(shiftedA_15__25_) );
  NOR2_X1 U2018 ( .A1(n160), .A2(n193), .ZN(shiftedA_15__24_) );
  NOR2_X1 U2019 ( .A1(n161), .A2(n193), .ZN(shiftedA_15__23_) );
  NOR2_X1 U2020 ( .A1(n162), .A2(n193), .ZN(shiftedA_15__22_) );
  NOR2_X1 U2021 ( .A1(n163), .A2(n193), .ZN(shiftedA_15__21_) );
  NOR2_X1 U2022 ( .A1(n164), .A2(n193), .ZN(shiftedA_15__20_) );
  NOR2_X1 U2023 ( .A1(n165), .A2(n193), .ZN(shiftedA_15__19_) );
  NOR2_X1 U2024 ( .A1(n166), .A2(n193), .ZN(shiftedA_15__18_) );
  NOR2_X1 U2025 ( .A1(n167), .A2(n193), .ZN(shiftedA_15__17_) );
  NOR2_X1 U2026 ( .A1(n168), .A2(n193), .ZN(shiftedA_15__16_) );
  NOR2_X1 U2027 ( .A1(n136), .A2(n193), .ZN(shiftedA_15__15_) );
  NOR2_X1 U2028 ( .A1(n139), .A2(n194), .ZN(shiftedA_14__44_) );
  NOR2_X1 U2029 ( .A1(n140), .A2(n194), .ZN(shiftedA_14__43_) );
  NOR2_X1 U2030 ( .A1(n141), .A2(n194), .ZN(shiftedA_14__42_) );
  NOR2_X1 U2031 ( .A1(n142), .A2(n194), .ZN(shiftedA_14__41_) );
  NOR2_X1 U2032 ( .A1(n143), .A2(n194), .ZN(shiftedA_14__40_) );
  NOR2_X1 U2033 ( .A1(n144), .A2(n194), .ZN(shiftedA_14__39_) );
  NOR2_X1 U2034 ( .A1(n145), .A2(n194), .ZN(shiftedA_14__38_) );
  NOR2_X1 U2035 ( .A1(n146), .A2(n194), .ZN(shiftedA_14__37_) );
  NOR2_X1 U2036 ( .A1(n147), .A2(n194), .ZN(shiftedA_14__36_) );
  NOR2_X1 U2037 ( .A1(n148), .A2(n194), .ZN(shiftedA_14__35_) );
  NOR2_X1 U2038 ( .A1(n149), .A2(n194), .ZN(shiftedA_14__34_) );
  NOR2_X1 U2039 ( .A1(n150), .A2(n194), .ZN(shiftedA_14__33_) );
  NOR2_X1 U2040 ( .A1(n151), .A2(n194), .ZN(shiftedA_14__32_) );
  NOR2_X1 U2041 ( .A1(n152), .A2(n194), .ZN(shiftedA_14__31_) );
  NOR2_X1 U2042 ( .A1(n153), .A2(n194), .ZN(shiftedA_14__30_) );
  NOR2_X1 U2043 ( .A1(n154), .A2(n194), .ZN(shiftedA_14__29_) );
  NOR2_X1 U2044 ( .A1(n155), .A2(n194), .ZN(shiftedA_14__28_) );
  NOR2_X1 U2045 ( .A1(n156), .A2(n194), .ZN(shiftedA_14__27_) );
  NOR2_X1 U2046 ( .A1(n157), .A2(n194), .ZN(shiftedA_14__26_) );
  NOR2_X1 U2047 ( .A1(n158), .A2(n194), .ZN(shiftedA_14__25_) );
  NOR2_X1 U2048 ( .A1(n159), .A2(n194), .ZN(shiftedA_14__24_) );
  NOR2_X1 U2049 ( .A1(n160), .A2(n194), .ZN(shiftedA_14__23_) );
  NOR2_X1 U2050 ( .A1(n161), .A2(n194), .ZN(shiftedA_14__22_) );
  NOR2_X1 U2051 ( .A1(n162), .A2(n194), .ZN(shiftedA_14__21_) );
  NOR2_X1 U2052 ( .A1(n163), .A2(n194), .ZN(shiftedA_14__20_) );
  NOR2_X1 U2053 ( .A1(n164), .A2(n194), .ZN(shiftedA_14__19_) );
  NOR2_X1 U2054 ( .A1(n165), .A2(n194), .ZN(shiftedA_14__18_) );
  NOR2_X1 U2055 ( .A1(n166), .A2(n194), .ZN(shiftedA_14__17_) );
  NOR2_X1 U2056 ( .A1(n167), .A2(n194), .ZN(shiftedA_14__16_) );
  NOR2_X1 U2057 ( .A1(n168), .A2(n194), .ZN(shiftedA_14__15_) );
  NOR2_X1 U2058 ( .A1(n136), .A2(n194), .ZN(shiftedA_14__14_) );
  NOR2_X1 U2059 ( .A1(n139), .A2(n195), .ZN(shiftedA_13__43_) );
  NOR2_X1 U2060 ( .A1(n140), .A2(n195), .ZN(shiftedA_13__42_) );
  NOR2_X1 U2061 ( .A1(n141), .A2(n195), .ZN(shiftedA_13__41_) );
  NOR2_X1 U2062 ( .A1(n142), .A2(n195), .ZN(shiftedA_13__40_) );
  NOR2_X1 U2063 ( .A1(n143), .A2(n195), .ZN(shiftedA_13__39_) );
  NOR2_X1 U2064 ( .A1(n144), .A2(n195), .ZN(shiftedA_13__38_) );
  NOR2_X1 U2065 ( .A1(n145), .A2(n195), .ZN(shiftedA_13__37_) );
  NOR2_X1 U2066 ( .A1(n146), .A2(n195), .ZN(shiftedA_13__36_) );
  NOR2_X1 U2067 ( .A1(n147), .A2(n195), .ZN(shiftedA_13__35_) );
  NOR2_X1 U2068 ( .A1(n148), .A2(n195), .ZN(shiftedA_13__34_) );
  NOR2_X1 U2069 ( .A1(n149), .A2(n195), .ZN(shiftedA_13__33_) );
  NOR2_X1 U2070 ( .A1(n150), .A2(n195), .ZN(shiftedA_13__32_) );
  NOR2_X1 U2071 ( .A1(n151), .A2(n195), .ZN(shiftedA_13__31_) );
  NOR2_X1 U2072 ( .A1(n152), .A2(n195), .ZN(shiftedA_13__30_) );
  NOR2_X1 U2073 ( .A1(n153), .A2(n195), .ZN(shiftedA_13__29_) );
  NOR2_X1 U2074 ( .A1(n154), .A2(n195), .ZN(shiftedA_13__28_) );
  NOR2_X1 U2075 ( .A1(n155), .A2(n195), .ZN(shiftedA_13__27_) );
  NOR2_X1 U2076 ( .A1(n156), .A2(n195), .ZN(shiftedA_13__26_) );
  NOR2_X1 U2077 ( .A1(n157), .A2(n195), .ZN(shiftedA_13__25_) );
  NOR2_X1 U2078 ( .A1(n158), .A2(n195), .ZN(shiftedA_13__24_) );
  NOR2_X1 U2079 ( .A1(n159), .A2(n195), .ZN(shiftedA_13__23_) );
  NOR2_X1 U2080 ( .A1(n160), .A2(n195), .ZN(shiftedA_13__22_) );
  NOR2_X1 U2081 ( .A1(n161), .A2(n195), .ZN(shiftedA_13__21_) );
  NOR2_X1 U2082 ( .A1(n162), .A2(n195), .ZN(shiftedA_13__20_) );
  NOR2_X1 U2083 ( .A1(n163), .A2(n195), .ZN(shiftedA_13__19_) );
  NOR2_X1 U2084 ( .A1(n164), .A2(n195), .ZN(shiftedA_13__18_) );
  NOR2_X1 U2085 ( .A1(n165), .A2(n195), .ZN(shiftedA_13__17_) );
  NOR2_X1 U2086 ( .A1(n166), .A2(n195), .ZN(shiftedA_13__16_) );
  NOR2_X1 U2087 ( .A1(n167), .A2(n195), .ZN(shiftedA_13__15_) );
  NOR2_X1 U2088 ( .A1(n168), .A2(n195), .ZN(shiftedA_13__14_) );
  NOR2_X1 U2089 ( .A1(n136), .A2(n195), .ZN(shiftedA_13__13_) );
  NOR2_X1 U2090 ( .A1(n139), .A2(n196), .ZN(shiftedA_12__42_) );
  NOR2_X1 U2091 ( .A1(n140), .A2(n196), .ZN(shiftedA_12__41_) );
  NOR2_X1 U2092 ( .A1(n141), .A2(n196), .ZN(shiftedA_12__40_) );
  NOR2_X1 U2093 ( .A1(n142), .A2(n196), .ZN(shiftedA_12__39_) );
  NOR2_X1 U2094 ( .A1(n143), .A2(n196), .ZN(shiftedA_12__38_) );
  NOR2_X1 U2095 ( .A1(n144), .A2(n196), .ZN(shiftedA_12__37_) );
  NOR2_X1 U2096 ( .A1(n145), .A2(n196), .ZN(shiftedA_12__36_) );
  NOR2_X1 U2097 ( .A1(n146), .A2(n196), .ZN(shiftedA_12__35_) );
  NOR2_X1 U2098 ( .A1(n147), .A2(n196), .ZN(shiftedA_12__34_) );
  NOR2_X1 U2099 ( .A1(n148), .A2(n196), .ZN(shiftedA_12__33_) );
  NOR2_X1 U2100 ( .A1(n149), .A2(n196), .ZN(shiftedA_12__32_) );
  NOR2_X1 U2101 ( .A1(n150), .A2(n196), .ZN(shiftedA_12__31_) );
  NOR2_X1 U2102 ( .A1(n151), .A2(n196), .ZN(shiftedA_12__30_) );
  NOR2_X1 U2103 ( .A1(n152), .A2(n196), .ZN(shiftedA_12__29_) );
  NOR2_X1 U2104 ( .A1(n153), .A2(n196), .ZN(shiftedA_12__28_) );
  NOR2_X1 U2105 ( .A1(n154), .A2(n196), .ZN(shiftedA_12__27_) );
  NOR2_X1 U2106 ( .A1(n155), .A2(n196), .ZN(shiftedA_12__26_) );
  NOR2_X1 U2107 ( .A1(n156), .A2(n196), .ZN(shiftedA_12__25_) );
  NOR2_X1 U2108 ( .A1(n157), .A2(n196), .ZN(shiftedA_12__24_) );
  NOR2_X1 U2109 ( .A1(n158), .A2(n196), .ZN(shiftedA_12__23_) );
  NOR2_X1 U2110 ( .A1(n159), .A2(n196), .ZN(shiftedA_12__22_) );
  NOR2_X1 U2111 ( .A1(n160), .A2(n196), .ZN(shiftedA_12__21_) );
  NOR2_X1 U2112 ( .A1(n161), .A2(n196), .ZN(shiftedA_12__20_) );
  NOR2_X1 U2113 ( .A1(n162), .A2(n196), .ZN(shiftedA_12__19_) );
  NOR2_X1 U2114 ( .A1(n163), .A2(n196), .ZN(shiftedA_12__18_) );
  NOR2_X1 U2115 ( .A1(n164), .A2(n196), .ZN(shiftedA_12__17_) );
  NOR2_X1 U2116 ( .A1(n165), .A2(n196), .ZN(shiftedA_12__16_) );
  NOR2_X1 U2117 ( .A1(n166), .A2(n196), .ZN(shiftedA_12__15_) );
  NOR2_X1 U2118 ( .A1(n167), .A2(n196), .ZN(shiftedA_12__14_) );
  NOR2_X1 U2119 ( .A1(n168), .A2(n196), .ZN(shiftedA_12__13_) );
  NOR2_X1 U2120 ( .A1(n136), .A2(n196), .ZN(shiftedA_12__12_) );
  NOR2_X1 U2121 ( .A1(n139), .A2(n197), .ZN(shiftedA_11__41_) );
  NOR2_X1 U2122 ( .A1(n140), .A2(n197), .ZN(shiftedA_11__40_) );
  NOR2_X1 U2123 ( .A1(n141), .A2(n197), .ZN(shiftedA_11__39_) );
  NOR2_X1 U2124 ( .A1(n142), .A2(n197), .ZN(shiftedA_11__38_) );
  NOR2_X1 U2125 ( .A1(n143), .A2(n197), .ZN(shiftedA_11__37_) );
  NOR2_X1 U2126 ( .A1(n144), .A2(n197), .ZN(shiftedA_11__36_) );
  NOR2_X1 U2127 ( .A1(n145), .A2(n197), .ZN(shiftedA_11__35_) );
  NOR2_X1 U2128 ( .A1(n146), .A2(n197), .ZN(shiftedA_11__34_) );
  NOR2_X1 U2129 ( .A1(n147), .A2(n197), .ZN(shiftedA_11__33_) );
  NOR2_X1 U2130 ( .A1(n148), .A2(n197), .ZN(shiftedA_11__32_) );
  NOR2_X1 U2131 ( .A1(n149), .A2(n197), .ZN(shiftedA_11__31_) );
  NOR2_X1 U2132 ( .A1(n150), .A2(n197), .ZN(shiftedA_11__30_) );
  NOR2_X1 U2133 ( .A1(n151), .A2(n197), .ZN(shiftedA_11__29_) );
  NOR2_X1 U2134 ( .A1(n152), .A2(n197), .ZN(shiftedA_11__28_) );
  NOR2_X1 U2135 ( .A1(n153), .A2(n197), .ZN(shiftedA_11__27_) );
  NOR2_X1 U2136 ( .A1(n154), .A2(n197), .ZN(shiftedA_11__26_) );
  NOR2_X1 U2137 ( .A1(n155), .A2(n197), .ZN(shiftedA_11__25_) );
  NOR2_X1 U2138 ( .A1(n156), .A2(n197), .ZN(shiftedA_11__24_) );
  NOR2_X1 U2139 ( .A1(n157), .A2(n197), .ZN(shiftedA_11__23_) );
  NOR2_X1 U2140 ( .A1(n158), .A2(n197), .ZN(shiftedA_11__22_) );
  NOR2_X1 U2141 ( .A1(n159), .A2(n197), .ZN(shiftedA_11__21_) );
  NOR2_X1 U2142 ( .A1(n160), .A2(n197), .ZN(shiftedA_11__20_) );
  NOR2_X1 U2143 ( .A1(n161), .A2(n197), .ZN(shiftedA_11__19_) );
  NOR2_X1 U2144 ( .A1(n162), .A2(n197), .ZN(shiftedA_11__18_) );
  NOR2_X1 U2145 ( .A1(n163), .A2(n197), .ZN(shiftedA_11__17_) );
  NOR2_X1 U2146 ( .A1(n164), .A2(n197), .ZN(shiftedA_11__16_) );
  NOR2_X1 U2147 ( .A1(n165), .A2(n197), .ZN(shiftedA_11__15_) );
  NOR2_X1 U2148 ( .A1(n166), .A2(n197), .ZN(shiftedA_11__14_) );
  NOR2_X1 U2149 ( .A1(n167), .A2(n197), .ZN(shiftedA_11__13_) );
  NOR2_X1 U2150 ( .A1(n168), .A2(n197), .ZN(shiftedA_11__12_) );
  NOR2_X1 U2151 ( .A1(n136), .A2(n197), .ZN(shiftedA_11__11_) );
  NOR2_X1 U2152 ( .A1(n139), .A2(n198), .ZN(shiftedA_10__40_) );
  NOR2_X1 U2153 ( .A1(n140), .A2(n198), .ZN(shiftedA_10__39_) );
  NOR2_X1 U2154 ( .A1(n141), .A2(n198), .ZN(shiftedA_10__38_) );
  NOR2_X1 U2155 ( .A1(n142), .A2(n198), .ZN(shiftedA_10__37_) );
  NOR2_X1 U2156 ( .A1(n143), .A2(n198), .ZN(shiftedA_10__36_) );
  NOR2_X1 U2157 ( .A1(n144), .A2(n198), .ZN(shiftedA_10__35_) );
  NOR2_X1 U2158 ( .A1(n145), .A2(n198), .ZN(shiftedA_10__34_) );
  NOR2_X1 U2159 ( .A1(n146), .A2(n198), .ZN(shiftedA_10__33_) );
  NOR2_X1 U2160 ( .A1(n147), .A2(n198), .ZN(shiftedA_10__32_) );
  NOR2_X1 U2161 ( .A1(n148), .A2(n198), .ZN(shiftedA_10__31_) );
  NOR2_X1 U2162 ( .A1(n149), .A2(n198), .ZN(shiftedA_10__30_) );
  NOR2_X1 U2163 ( .A1(n150), .A2(n198), .ZN(shiftedA_10__29_) );
  NOR2_X1 U2164 ( .A1(n151), .A2(n198), .ZN(shiftedA_10__28_) );
  NOR2_X1 U2165 ( .A1(n152), .A2(n198), .ZN(shiftedA_10__27_) );
  NOR2_X1 U2166 ( .A1(n153), .A2(n198), .ZN(shiftedA_10__26_) );
  NOR2_X1 U2167 ( .A1(n154), .A2(n198), .ZN(shiftedA_10__25_) );
  NOR2_X1 U2168 ( .A1(n155), .A2(n198), .ZN(shiftedA_10__24_) );
  NOR2_X1 U2169 ( .A1(n156), .A2(n198), .ZN(shiftedA_10__23_) );
  NOR2_X1 U2170 ( .A1(n157), .A2(n198), .ZN(shiftedA_10__22_) );
  NOR2_X1 U2171 ( .A1(n158), .A2(n198), .ZN(shiftedA_10__21_) );
  NOR2_X1 U2172 ( .A1(n159), .A2(n198), .ZN(shiftedA_10__20_) );
  NOR2_X1 U2173 ( .A1(n160), .A2(n198), .ZN(shiftedA_10__19_) );
  NOR2_X1 U2174 ( .A1(n161), .A2(n198), .ZN(shiftedA_10__18_) );
  NOR2_X1 U2175 ( .A1(n162), .A2(n198), .ZN(shiftedA_10__17_) );
  NOR2_X1 U2176 ( .A1(n163), .A2(n198), .ZN(shiftedA_10__16_) );
  NOR2_X1 U2177 ( .A1(n164), .A2(n198), .ZN(shiftedA_10__15_) );
  NOR2_X1 U2178 ( .A1(n165), .A2(n198), .ZN(shiftedA_10__14_) );
  NOR2_X1 U2179 ( .A1(n166), .A2(n198), .ZN(shiftedA_10__13_) );
  NOR2_X1 U2180 ( .A1(n167), .A2(n198), .ZN(shiftedA_10__12_) );
  NOR2_X1 U2181 ( .A1(n168), .A2(n198), .ZN(shiftedA_10__11_) );
  NOR2_X1 U2182 ( .A1(n136), .A2(n198), .ZN(shiftedA_10__10_) );
  NOR2_X1 U2183 ( .A1(n160), .A2(n199), .ZN(shiftedA_0__9_) );
  NOR2_X1 U2184 ( .A1(n161), .A2(n199), .ZN(shiftedA_0__8_) );
  NOR2_X1 U2185 ( .A1(n162), .A2(n199), .ZN(shiftedA_0__7_) );
  NOR2_X1 U2186 ( .A1(n163), .A2(n199), .ZN(shiftedA_0__6_) );
  NOR2_X1 U2187 ( .A1(n164), .A2(n199), .ZN(shiftedA_0__5_) );
  NOR2_X1 U2188 ( .A1(n165), .A2(n199), .ZN(shiftedA_0__4_) );
  NOR2_X1 U2189 ( .A1(n166), .A2(n199), .ZN(shiftedA_0__3_) );
  NOR2_X1 U2190 ( .A1(n139), .A2(n199), .ZN(shiftedA_0__30_) );
  NOR2_X1 U2191 ( .A1(n167), .A2(n199), .ZN(shiftedA_0__2_) );
  NOR2_X1 U2192 ( .A1(n140), .A2(n199), .ZN(shiftedA_0__29_) );
  NOR2_X1 U2193 ( .A1(n141), .A2(n199), .ZN(shiftedA_0__28_) );
  NOR2_X1 U2194 ( .A1(n142), .A2(n199), .ZN(shiftedA_0__27_) );
  NOR2_X1 U2195 ( .A1(n143), .A2(n199), .ZN(shiftedA_0__26_) );
  NOR2_X1 U2196 ( .A1(n144), .A2(n199), .ZN(shiftedA_0__25_) );
  NOR2_X1 U2197 ( .A1(n145), .A2(n199), .ZN(shiftedA_0__24_) );
  NOR2_X1 U2198 ( .A1(n146), .A2(n199), .ZN(shiftedA_0__23_) );
  NOR2_X1 U2199 ( .A1(n147), .A2(n199), .ZN(shiftedA_0__22_) );
  NOR2_X1 U2200 ( .A1(n148), .A2(n199), .ZN(shiftedA_0__21_) );
  NOR2_X1 U2201 ( .A1(n149), .A2(n199), .ZN(shiftedA_0__20_) );
  NOR2_X1 U2202 ( .A1(n168), .A2(n199), .ZN(shiftedA_0__1_) );
  NOR2_X1 U2203 ( .A1(n150), .A2(n199), .ZN(shiftedA_0__19_) );
  NOR2_X1 U2204 ( .A1(n151), .A2(n199), .ZN(shiftedA_0__18_) );
  NOR2_X1 U2205 ( .A1(n152), .A2(n199), .ZN(shiftedA_0__17_) );
  NOR2_X1 U2206 ( .A1(n153), .A2(n199), .ZN(shiftedA_0__16_) );
  NOR2_X1 U2207 ( .A1(n154), .A2(n199), .ZN(shiftedA_0__15_) );
  NOR2_X1 U2208 ( .A1(n155), .A2(n199), .ZN(shiftedA_0__14_) );
  NOR2_X1 U2209 ( .A1(n156), .A2(n199), .ZN(shiftedA_0__13_) );
  NOR2_X1 U2210 ( .A1(n157), .A2(n199), .ZN(shiftedA_0__12_) );
  NOR2_X1 U2211 ( .A1(n158), .A2(n199), .ZN(shiftedA_0__11_) );
  NOR2_X1 U2212 ( .A1(n159), .A2(n199), .ZN(shiftedA_0__10_) );
  NOR2_X1 U2213 ( .A1(n136), .A2(n199), .ZN(shiftedA_0__0_) );
endmodule


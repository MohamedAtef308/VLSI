
module FullAdder_0 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_1 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_2 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_3 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_4 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_5 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_6 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_7 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_8 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_9 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_10 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_11 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_12 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_13 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_14 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_15 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_16 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_17 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_18 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_19 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_20 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_21 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_22 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_23 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_24 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_25 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_26 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_27 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_28 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_29 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_30 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_31 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_32 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_33 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_34 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_35 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_36 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_37 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_38 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_39 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_40 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_41 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_42 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_43 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_44 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_45 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_46 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_47 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_48 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_49 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_50 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_51 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_52 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_53 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_54 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_55 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_56 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_57 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_58 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_59 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_60 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_61 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_62 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module FullAdder_63 ( a, b, cin, sum, cout );
  input a, b, cin;
  output sum, cout;
  wire   n1, n2;

  XOR2_X1 U1 ( .A(cin), .B(n1), .Z(sum) );
  INV_X1 U2 ( .A(n2), .ZN(cout) );
  AOI22_X1 U3 ( .A1(b), .A2(a), .B1(n1), .B2(cin), .ZN(n2) );
  XOR2_X1 U4 ( .A(a), .B(b), .Z(n1) );
endmodule


module CRAdder_64 ( a, b, cin, sum, cout, overflow );
  input [63:0] a;
  input [63:0] b;
  output [63:0] sum;
  input cin;
  output cout, overflow;
  wire   n3, n4;
  wire   [62:0] passCout;

  FullAdder_0 bit0 ( .a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(
        passCout[0]) );
  FullAdder_63 bit_gen_1__bit ( .a(a[1]), .b(b[1]), .cin(passCout[0]), .sum(
        sum[1]), .cout(passCout[1]) );
  FullAdder_62 bit_gen_2__bit ( .a(a[2]), .b(b[2]), .cin(passCout[1]), .sum(
        sum[2]), .cout(passCout[2]) );
  FullAdder_61 bit_gen_3__bit ( .a(a[3]), .b(b[3]), .cin(passCout[2]), .sum(
        sum[3]), .cout(passCout[3]) );
  FullAdder_60 bit_gen_4__bit ( .a(a[4]), .b(b[4]), .cin(passCout[3]), .sum(
        sum[4]), .cout(passCout[4]) );
  FullAdder_59 bit_gen_5__bit ( .a(a[5]), .b(b[5]), .cin(passCout[4]), .sum(
        sum[5]), .cout(passCout[5]) );
  FullAdder_58 bit_gen_6__bit ( .a(a[6]), .b(b[6]), .cin(passCout[5]), .sum(
        sum[6]), .cout(passCout[6]) );
  FullAdder_57 bit_gen_7__bit ( .a(a[7]), .b(b[7]), .cin(passCout[6]), .sum(
        sum[7]), .cout(passCout[7]) );
  FullAdder_56 bit_gen_8__bit ( .a(a[8]), .b(b[8]), .cin(passCout[7]), .sum(
        sum[8]), .cout(passCout[8]) );
  FullAdder_55 bit_gen_9__bit ( .a(a[9]), .b(b[9]), .cin(passCout[8]), .sum(
        sum[9]), .cout(passCout[9]) );
  FullAdder_54 bit_gen_10__bit ( .a(a[10]), .b(b[10]), .cin(passCout[9]), 
        .sum(sum[10]), .cout(passCout[10]) );
  FullAdder_53 bit_gen_11__bit ( .a(a[11]), .b(b[11]), .cin(passCout[10]), 
        .sum(sum[11]), .cout(passCout[11]) );
  FullAdder_52 bit_gen_12__bit ( .a(a[12]), .b(b[12]), .cin(passCout[11]), 
        .sum(sum[12]), .cout(passCout[12]) );
  FullAdder_51 bit_gen_13__bit ( .a(a[13]), .b(b[13]), .cin(passCout[12]), 
        .sum(sum[13]), .cout(passCout[13]) );
  FullAdder_50 bit_gen_14__bit ( .a(a[14]), .b(b[14]), .cin(passCout[13]), 
        .sum(sum[14]), .cout(passCout[14]) );
  FullAdder_49 bit_gen_15__bit ( .a(a[15]), .b(b[15]), .cin(passCout[14]), 
        .sum(sum[15]), .cout(passCout[15]) );
  FullAdder_48 bit_gen_16__bit ( .a(a[16]), .b(b[16]), .cin(passCout[15]), 
        .sum(sum[16]), .cout(passCout[16]) );
  FullAdder_47 bit_gen_17__bit ( .a(a[17]), .b(b[17]), .cin(passCout[16]), 
        .sum(sum[17]), .cout(passCout[17]) );
  FullAdder_46 bit_gen_18__bit ( .a(a[18]), .b(b[18]), .cin(passCout[17]), 
        .sum(sum[18]), .cout(passCout[18]) );
  FullAdder_45 bit_gen_19__bit ( .a(a[19]), .b(b[19]), .cin(passCout[18]), 
        .sum(sum[19]), .cout(passCout[19]) );
  FullAdder_44 bit_gen_20__bit ( .a(a[20]), .b(b[20]), .cin(passCout[19]), 
        .sum(sum[20]), .cout(passCout[20]) );
  FullAdder_43 bit_gen_21__bit ( .a(a[21]), .b(b[21]), .cin(passCout[20]), 
        .sum(sum[21]), .cout(passCout[21]) );
  FullAdder_42 bit_gen_22__bit ( .a(a[22]), .b(b[22]), .cin(passCout[21]), 
        .sum(sum[22]), .cout(passCout[22]) );
  FullAdder_41 bit_gen_23__bit ( .a(a[23]), .b(b[23]), .cin(passCout[22]), 
        .sum(sum[23]), .cout(passCout[23]) );
  FullAdder_40 bit_gen_24__bit ( .a(a[24]), .b(b[24]), .cin(passCout[23]), 
        .sum(sum[24]), .cout(passCout[24]) );
  FullAdder_39 bit_gen_25__bit ( .a(a[25]), .b(b[25]), .cin(passCout[24]), 
        .sum(sum[25]), .cout(passCout[25]) );
  FullAdder_38 bit_gen_26__bit ( .a(a[26]), .b(b[26]), .cin(passCout[25]), 
        .sum(sum[26]), .cout(passCout[26]) );
  FullAdder_37 bit_gen_27__bit ( .a(a[27]), .b(b[27]), .cin(passCout[26]), 
        .sum(sum[27]), .cout(passCout[27]) );
  FullAdder_36 bit_gen_28__bit ( .a(a[28]), .b(b[28]), .cin(passCout[27]), 
        .sum(sum[28]), .cout(passCout[28]) );
  FullAdder_35 bit_gen_29__bit ( .a(a[29]), .b(b[29]), .cin(passCout[28]), 
        .sum(sum[29]), .cout(passCout[29]) );
  FullAdder_34 bit_gen_30__bit ( .a(a[30]), .b(b[30]), .cin(passCout[29]), 
        .sum(sum[30]), .cout(passCout[30]) );
  FullAdder_33 bit_gen_31__bit ( .a(a[31]), .b(b[31]), .cin(passCout[30]), 
        .sum(sum[31]), .cout(passCout[31]) );
  FullAdder_32 bit_gen_32__bit ( .a(a[32]), .b(b[32]), .cin(passCout[31]), 
        .sum(sum[32]), .cout(passCout[32]) );
  FullAdder_31 bit_gen_33__bit ( .a(a[33]), .b(b[33]), .cin(passCout[32]), 
        .sum(sum[33]), .cout(passCout[33]) );
  FullAdder_30 bit_gen_34__bit ( .a(a[34]), .b(b[34]), .cin(passCout[33]), 
        .sum(sum[34]), .cout(passCout[34]) );
  FullAdder_29 bit_gen_35__bit ( .a(a[35]), .b(b[35]), .cin(passCout[34]), 
        .sum(sum[35]), .cout(passCout[35]) );
  FullAdder_28 bit_gen_36__bit ( .a(a[36]), .b(b[36]), .cin(passCout[35]), 
        .sum(sum[36]), .cout(passCout[36]) );
  FullAdder_27 bit_gen_37__bit ( .a(a[37]), .b(b[37]), .cin(passCout[36]), 
        .sum(sum[37]), .cout(passCout[37]) );
  FullAdder_26 bit_gen_38__bit ( .a(a[38]), .b(b[38]), .cin(passCout[37]), 
        .sum(sum[38]), .cout(passCout[38]) );
  FullAdder_25 bit_gen_39__bit ( .a(a[39]), .b(b[39]), .cin(passCout[38]), 
        .sum(sum[39]), .cout(passCout[39]) );
  FullAdder_24 bit_gen_40__bit ( .a(a[40]), .b(b[40]), .cin(passCout[39]), 
        .sum(sum[40]), .cout(passCout[40]) );
  FullAdder_23 bit_gen_41__bit ( .a(a[41]), .b(b[41]), .cin(passCout[40]), 
        .sum(sum[41]), .cout(passCout[41]) );
  FullAdder_22 bit_gen_42__bit ( .a(a[42]), .b(b[42]), .cin(passCout[41]), 
        .sum(sum[42]), .cout(passCout[42]) );
  FullAdder_21 bit_gen_43__bit ( .a(a[43]), .b(b[43]), .cin(passCout[42]), 
        .sum(sum[43]), .cout(passCout[43]) );
  FullAdder_20 bit_gen_44__bit ( .a(a[44]), .b(b[44]), .cin(passCout[43]), 
        .sum(sum[44]), .cout(passCout[44]) );
  FullAdder_19 bit_gen_45__bit ( .a(a[45]), .b(b[45]), .cin(passCout[44]), 
        .sum(sum[45]), .cout(passCout[45]) );
  FullAdder_18 bit_gen_46__bit ( .a(a[46]), .b(b[46]), .cin(passCout[45]), 
        .sum(sum[46]), .cout(passCout[46]) );
  FullAdder_17 bit_gen_47__bit ( .a(a[47]), .b(b[47]), .cin(passCout[46]), 
        .sum(sum[47]), .cout(passCout[47]) );
  FullAdder_16 bit_gen_48__bit ( .a(a[48]), .b(b[48]), .cin(passCout[47]), 
        .sum(sum[48]), .cout(passCout[48]) );
  FullAdder_15 bit_gen_49__bit ( .a(a[49]), .b(b[49]), .cin(passCout[48]), 
        .sum(sum[49]), .cout(passCout[49]) );
  FullAdder_14 bit_gen_50__bit ( .a(a[50]), .b(b[50]), .cin(passCout[49]), 
        .sum(sum[50]), .cout(passCout[50]) );
  FullAdder_13 bit_gen_51__bit ( .a(a[51]), .b(b[51]), .cin(passCout[50]), 
        .sum(sum[51]), .cout(passCout[51]) );
  FullAdder_12 bit_gen_52__bit ( .a(a[52]), .b(b[52]), .cin(passCout[51]), 
        .sum(sum[52]), .cout(passCout[52]) );
  FullAdder_11 bit_gen_53__bit ( .a(a[53]), .b(b[53]), .cin(passCout[52]), 
        .sum(sum[53]), .cout(passCout[53]) );
  FullAdder_10 bit_gen_54__bit ( .a(a[54]), .b(b[54]), .cin(passCout[53]), 
        .sum(sum[54]), .cout(passCout[54]) );
  FullAdder_9 bit_gen_55__bit ( .a(a[55]), .b(b[55]), .cin(passCout[54]), 
        .sum(sum[55]), .cout(passCout[55]) );
  FullAdder_8 bit_gen_56__bit ( .a(a[56]), .b(b[56]), .cin(passCout[55]), 
        .sum(sum[56]), .cout(passCout[56]) );
  FullAdder_7 bit_gen_57__bit ( .a(a[57]), .b(b[57]), .cin(passCout[56]), 
        .sum(sum[57]), .cout(passCout[57]) );
  FullAdder_6 bit_gen_58__bit ( .a(a[58]), .b(b[58]), .cin(passCout[57]), 
        .sum(sum[58]), .cout(passCout[58]) );
  FullAdder_5 bit_gen_59__bit ( .a(a[59]), .b(b[59]), .cin(passCout[58]), 
        .sum(sum[59]), .cout(passCout[59]) );
  FullAdder_4 bit_gen_60__bit ( .a(a[60]), .b(b[60]), .cin(passCout[59]), 
        .sum(sum[60]), .cout(passCout[60]) );
  FullAdder_3 bit_gen_61__bit ( .a(a[61]), .b(b[61]), .cin(passCout[60]), 
        .sum(sum[61]), .cout(passCout[61]) );
  FullAdder_2 bit_gen_62__bit ( .a(a[62]), .b(b[62]), .cin(passCout[61]), 
        .sum(sum[62]), .cout(passCout[62]) );
  FullAdder_1 bit63 ( .a(a[63]), .b(b[63]), .cin(passCout[62]), .sum(sum[63]), 
        .cout(cout) );
  NOR2_X1 U4 ( .A1(n3), .A2(n4), .ZN(overflow) );
  XOR2_X1 U5 ( .A(b[63]), .B(a[63]), .Z(n4) );
  XNOR2_X1 U6 ( .A(a[63]), .B(sum[63]), .ZN(n3) );
endmodule

